
module dummy_top(output dum_out);

//wire dum_out;


wire [6143:0] A,B;

assign dum_out=B[6000];

wire k;

coder_interleaver dummy_inst(
		.cin(A),
		.K_eq_6144(k),
		.cout(B)
	);
	
	
endmodule 