module mux6144(
arr,
in,
r
);

input [13:0] in;
input [6143:0] arr;

output r;


wire r1_1;
assign r1_1 = in[0]? arr[1] : arr[0];
wire r1_2;
assign r1_2 = in[0]? arr[3] : arr[2];
wire r1_3;
assign r1_3 = in[0]? arr[5] : arr[4];
wire r1_4;
assign r1_4 = in[0]? arr[7] : arr[6];
wire r1_5;
assign r1_5 = in[0]? arr[9] : arr[8];
wire r1_6;
assign r1_6 = in[0]? arr[11] : arr[10];
wire r1_7;
assign r1_7 = in[0]? arr[13] : arr[12];
wire r1_8;
assign r1_8 = in[0]? arr[15] : arr[14];
wire r1_9;
assign r1_9 = in[0]? arr[17] : arr[16];
wire r1_10;
assign r1_10 = in[0]? arr[19] : arr[18];
wire r1_11;
assign r1_11 = in[0]? arr[21] : arr[20];
wire r1_12;
assign r1_12 = in[0]? arr[23] : arr[22];
wire r1_13;
assign r1_13 = in[0]? arr[25] : arr[24];
wire r1_14;
assign r1_14 = in[0]? arr[27] : arr[26];
wire r1_15;
assign r1_15 = in[0]? arr[29] : arr[28];
wire r1_16;
assign r1_16 = in[0]? arr[31] : arr[30];
wire r1_17;
assign r1_17 = in[0]? arr[33] : arr[32];
wire r1_18;
assign r1_18 = in[0]? arr[35] : arr[34];
wire r1_19;
assign r1_19 = in[0]? arr[37] : arr[36];
wire r1_20;
assign r1_20 = in[0]? arr[39] : arr[38];
wire r1_21;
assign r1_21 = in[0]? arr[41] : arr[40];
wire r1_22;
assign r1_22 = in[0]? arr[43] : arr[42];
wire r1_23;
assign r1_23 = in[0]? arr[45] : arr[44];
wire r1_24;
assign r1_24 = in[0]? arr[47] : arr[46];
wire r1_25;
assign r1_25 = in[0]? arr[49] : arr[48];
wire r1_26;
assign r1_26 = in[0]? arr[51] : arr[50];
wire r1_27;
assign r1_27 = in[0]? arr[53] : arr[52];
wire r1_28;
assign r1_28 = in[0]? arr[55] : arr[54];
wire r1_29;
assign r1_29 = in[0]? arr[57] : arr[56];
wire r1_30;
assign r1_30 = in[0]? arr[59] : arr[58];
wire r1_31;
assign r1_31 = in[0]? arr[61] : arr[60];
wire r1_32;
assign r1_32 = in[0]? arr[63] : arr[62];
wire r1_33;
assign r1_33 = in[0]? arr[65] : arr[64];
wire r1_34;
assign r1_34 = in[0]? arr[67] : arr[66];
wire r1_35;
assign r1_35 = in[0]? arr[69] : arr[68];
wire r1_36;
assign r1_36 = in[0]? arr[71] : arr[70];
wire r1_37;
assign r1_37 = in[0]? arr[73] : arr[72];
wire r1_38;
assign r1_38 = in[0]? arr[75] : arr[74];
wire r1_39;
assign r1_39 = in[0]? arr[77] : arr[76];
wire r1_40;
assign r1_40 = in[0]? arr[79] : arr[78];
wire r1_41;
assign r1_41 = in[0]? arr[81] : arr[80];
wire r1_42;
assign r1_42 = in[0]? arr[83] : arr[82];
wire r1_43;
assign r1_43 = in[0]? arr[85] : arr[84];
wire r1_44;
assign r1_44 = in[0]? arr[87] : arr[86];
wire r1_45;
assign r1_45 = in[0]? arr[89] : arr[88];
wire r1_46;
assign r1_46 = in[0]? arr[91] : arr[90];
wire r1_47;
assign r1_47 = in[0]? arr[93] : arr[92];
wire r1_48;
assign r1_48 = in[0]? arr[95] : arr[94];
wire r1_49;
assign r1_49 = in[0]? arr[97] : arr[96];
wire r1_50;
assign r1_50 = in[0]? arr[99] : arr[98];
wire r1_51;
assign r1_51 = in[0]? arr[101] : arr[100];
wire r1_52;
assign r1_52 = in[0]? arr[103] : arr[102];
wire r1_53;
assign r1_53 = in[0]? arr[105] : arr[104];
wire r1_54;
assign r1_54 = in[0]? arr[107] : arr[106];
wire r1_55;
assign r1_55 = in[0]? arr[109] : arr[108];
wire r1_56;
assign r1_56 = in[0]? arr[111] : arr[110];
wire r1_57;
assign r1_57 = in[0]? arr[113] : arr[112];
wire r1_58;
assign r1_58 = in[0]? arr[115] : arr[114];
wire r1_59;
assign r1_59 = in[0]? arr[117] : arr[116];
wire r1_60;
assign r1_60 = in[0]? arr[119] : arr[118];
wire r1_61;
assign r1_61 = in[0]? arr[121] : arr[120];
wire r1_62;
assign r1_62 = in[0]? arr[123] : arr[122];
wire r1_63;
assign r1_63 = in[0]? arr[125] : arr[124];
wire r1_64;
assign r1_64 = in[0]? arr[127] : arr[126];
wire r1_65;
assign r1_65 = in[0]? arr[129] : arr[128];
wire r1_66;
assign r1_66 = in[0]? arr[131] : arr[130];
wire r1_67;
assign r1_67 = in[0]? arr[133] : arr[132];
wire r1_68;
assign r1_68 = in[0]? arr[135] : arr[134];
wire r1_69;
assign r1_69 = in[0]? arr[137] : arr[136];
wire r1_70;
assign r1_70 = in[0]? arr[139] : arr[138];
wire r1_71;
assign r1_71 = in[0]? arr[141] : arr[140];
wire r1_72;
assign r1_72 = in[0]? arr[143] : arr[142];
wire r1_73;
assign r1_73 = in[0]? arr[145] : arr[144];
wire r1_74;
assign r1_74 = in[0]? arr[147] : arr[146];
wire r1_75;
assign r1_75 = in[0]? arr[149] : arr[148];
wire r1_76;
assign r1_76 = in[0]? arr[151] : arr[150];
wire r1_77;
assign r1_77 = in[0]? arr[153] : arr[152];
wire r1_78;
assign r1_78 = in[0]? arr[155] : arr[154];
wire r1_79;
assign r1_79 = in[0]? arr[157] : arr[156];
wire r1_80;
assign r1_80 = in[0]? arr[159] : arr[158];
wire r1_81;
assign r1_81 = in[0]? arr[161] : arr[160];
wire r1_82;
assign r1_82 = in[0]? arr[163] : arr[162];
wire r1_83;
assign r1_83 = in[0]? arr[165] : arr[164];
wire r1_84;
assign r1_84 = in[0]? arr[167] : arr[166];
wire r1_85;
assign r1_85 = in[0]? arr[169] : arr[168];
wire r1_86;
assign r1_86 = in[0]? arr[171] : arr[170];
wire r1_87;
assign r1_87 = in[0]? arr[173] : arr[172];
wire r1_88;
assign r1_88 = in[0]? arr[175] : arr[174];
wire r1_89;
assign r1_89 = in[0]? arr[177] : arr[176];
wire r1_90;
assign r1_90 = in[0]? arr[179] : arr[178];
wire r1_91;
assign r1_91 = in[0]? arr[181] : arr[180];
wire r1_92;
assign r1_92 = in[0]? arr[183] : arr[182];
wire r1_93;
assign r1_93 = in[0]? arr[185] : arr[184];
wire r1_94;
assign r1_94 = in[0]? arr[187] : arr[186];
wire r1_95;
assign r1_95 = in[0]? arr[189] : arr[188];
wire r1_96;
assign r1_96 = in[0]? arr[191] : arr[190];
wire r1_97;
assign r1_97 = in[0]? arr[193] : arr[192];
wire r1_98;
assign r1_98 = in[0]? arr[195] : arr[194];
wire r1_99;
assign r1_99 = in[0]? arr[197] : arr[196];
wire r1_100;
assign r1_100 = in[0]? arr[199] : arr[198];
wire r1_101;
assign r1_101 = in[0]? arr[201] : arr[200];
wire r1_102;
assign r1_102 = in[0]? arr[203] : arr[202];
wire r1_103;
assign r1_103 = in[0]? arr[205] : arr[204];
wire r1_104;
assign r1_104 = in[0]? arr[207] : arr[206];
wire r1_105;
assign r1_105 = in[0]? arr[209] : arr[208];
wire r1_106;
assign r1_106 = in[0]? arr[211] : arr[210];
wire r1_107;
assign r1_107 = in[0]? arr[213] : arr[212];
wire r1_108;
assign r1_108 = in[0]? arr[215] : arr[214];
wire r1_109;
assign r1_109 = in[0]? arr[217] : arr[216];
wire r1_110;
assign r1_110 = in[0]? arr[219] : arr[218];
wire r1_111;
assign r1_111 = in[0]? arr[221] : arr[220];
wire r1_112;
assign r1_112 = in[0]? arr[223] : arr[222];
wire r1_113;
assign r1_113 = in[0]? arr[225] : arr[224];
wire r1_114;
assign r1_114 = in[0]? arr[227] : arr[226];
wire r1_115;
assign r1_115 = in[0]? arr[229] : arr[228];
wire r1_116;
assign r1_116 = in[0]? arr[231] : arr[230];
wire r1_117;
assign r1_117 = in[0]? arr[233] : arr[232];
wire r1_118;
assign r1_118 = in[0]? arr[235] : arr[234];
wire r1_119;
assign r1_119 = in[0]? arr[237] : arr[236];
wire r1_120;
assign r1_120 = in[0]? arr[239] : arr[238];
wire r1_121;
assign r1_121 = in[0]? arr[241] : arr[240];
wire r1_122;
assign r1_122 = in[0]? arr[243] : arr[242];
wire r1_123;
assign r1_123 = in[0]? arr[245] : arr[244];
wire r1_124;
assign r1_124 = in[0]? arr[247] : arr[246];
wire r1_125;
assign r1_125 = in[0]? arr[249] : arr[248];
wire r1_126;
assign r1_126 = in[0]? arr[251] : arr[250];
wire r1_127;
assign r1_127 = in[0]? arr[253] : arr[252];
wire r1_128;
assign r1_128 = in[0]? arr[255] : arr[254];
wire r1_129;
assign r1_129 = in[0]? arr[257] : arr[256];
wire r1_130;
assign r1_130 = in[0]? arr[259] : arr[258];
wire r1_131;
assign r1_131 = in[0]? arr[261] : arr[260];
wire r1_132;
assign r1_132 = in[0]? arr[263] : arr[262];
wire r1_133;
assign r1_133 = in[0]? arr[265] : arr[264];
wire r1_134;
assign r1_134 = in[0]? arr[267] : arr[266];
wire r1_135;
assign r1_135 = in[0]? arr[269] : arr[268];
wire r1_136;
assign r1_136 = in[0]? arr[271] : arr[270];
wire r1_137;
assign r1_137 = in[0]? arr[273] : arr[272];
wire r1_138;
assign r1_138 = in[0]? arr[275] : arr[274];
wire r1_139;
assign r1_139 = in[0]? arr[277] : arr[276];
wire r1_140;
assign r1_140 = in[0]? arr[279] : arr[278];
wire r1_141;
assign r1_141 = in[0]? arr[281] : arr[280];
wire r1_142;
assign r1_142 = in[0]? arr[283] : arr[282];
wire r1_143;
assign r1_143 = in[0]? arr[285] : arr[284];
wire r1_144;
assign r1_144 = in[0]? arr[287] : arr[286];
wire r1_145;
assign r1_145 = in[0]? arr[289] : arr[288];
wire r1_146;
assign r1_146 = in[0]? arr[291] : arr[290];
wire r1_147;
assign r1_147 = in[0]? arr[293] : arr[292];
wire r1_148;
assign r1_148 = in[0]? arr[295] : arr[294];
wire r1_149;
assign r1_149 = in[0]? arr[297] : arr[296];
wire r1_150;
assign r1_150 = in[0]? arr[299] : arr[298];
wire r1_151;
assign r1_151 = in[0]? arr[301] : arr[300];
wire r1_152;
assign r1_152 = in[0]? arr[303] : arr[302];
wire r1_153;
assign r1_153 = in[0]? arr[305] : arr[304];
wire r1_154;
assign r1_154 = in[0]? arr[307] : arr[306];
wire r1_155;
assign r1_155 = in[0]? arr[309] : arr[308];
wire r1_156;
assign r1_156 = in[0]? arr[311] : arr[310];
wire r1_157;
assign r1_157 = in[0]? arr[313] : arr[312];
wire r1_158;
assign r1_158 = in[0]? arr[315] : arr[314];
wire r1_159;
assign r1_159 = in[0]? arr[317] : arr[316];
wire r1_160;
assign r1_160 = in[0]? arr[319] : arr[318];
wire r1_161;
assign r1_161 = in[0]? arr[321] : arr[320];
wire r1_162;
assign r1_162 = in[0]? arr[323] : arr[322];
wire r1_163;
assign r1_163 = in[0]? arr[325] : arr[324];
wire r1_164;
assign r1_164 = in[0]? arr[327] : arr[326];
wire r1_165;
assign r1_165 = in[0]? arr[329] : arr[328];
wire r1_166;
assign r1_166 = in[0]? arr[331] : arr[330];
wire r1_167;
assign r1_167 = in[0]? arr[333] : arr[332];
wire r1_168;
assign r1_168 = in[0]? arr[335] : arr[334];
wire r1_169;
assign r1_169 = in[0]? arr[337] : arr[336];
wire r1_170;
assign r1_170 = in[0]? arr[339] : arr[338];
wire r1_171;
assign r1_171 = in[0]? arr[341] : arr[340];
wire r1_172;
assign r1_172 = in[0]? arr[343] : arr[342];
wire r1_173;
assign r1_173 = in[0]? arr[345] : arr[344];
wire r1_174;
assign r1_174 = in[0]? arr[347] : arr[346];
wire r1_175;
assign r1_175 = in[0]? arr[349] : arr[348];
wire r1_176;
assign r1_176 = in[0]? arr[351] : arr[350];
wire r1_177;
assign r1_177 = in[0]? arr[353] : arr[352];
wire r1_178;
assign r1_178 = in[0]? arr[355] : arr[354];
wire r1_179;
assign r1_179 = in[0]? arr[357] : arr[356];
wire r1_180;
assign r1_180 = in[0]? arr[359] : arr[358];
wire r1_181;
assign r1_181 = in[0]? arr[361] : arr[360];
wire r1_182;
assign r1_182 = in[0]? arr[363] : arr[362];
wire r1_183;
assign r1_183 = in[0]? arr[365] : arr[364];
wire r1_184;
assign r1_184 = in[0]? arr[367] : arr[366];
wire r1_185;
assign r1_185 = in[0]? arr[369] : arr[368];
wire r1_186;
assign r1_186 = in[0]? arr[371] : arr[370];
wire r1_187;
assign r1_187 = in[0]? arr[373] : arr[372];
wire r1_188;
assign r1_188 = in[0]? arr[375] : arr[374];
wire r1_189;
assign r1_189 = in[0]? arr[377] : arr[376];
wire r1_190;
assign r1_190 = in[0]? arr[379] : arr[378];
wire r1_191;
assign r1_191 = in[0]? arr[381] : arr[380];
wire r1_192;
assign r1_192 = in[0]? arr[383] : arr[382];
wire r1_193;
assign r1_193 = in[0]? arr[385] : arr[384];
wire r1_194;
assign r1_194 = in[0]? arr[387] : arr[386];
wire r1_195;
assign r1_195 = in[0]? arr[389] : arr[388];
wire r1_196;
assign r1_196 = in[0]? arr[391] : arr[390];
wire r1_197;
assign r1_197 = in[0]? arr[393] : arr[392];
wire r1_198;
assign r1_198 = in[0]? arr[395] : arr[394];
wire r1_199;
assign r1_199 = in[0]? arr[397] : arr[396];
wire r1_200;
assign r1_200 = in[0]? arr[399] : arr[398];
wire r1_201;
assign r1_201 = in[0]? arr[401] : arr[400];
wire r1_202;
assign r1_202 = in[0]? arr[403] : arr[402];
wire r1_203;
assign r1_203 = in[0]? arr[405] : arr[404];
wire r1_204;
assign r1_204 = in[0]? arr[407] : arr[406];
wire r1_205;
assign r1_205 = in[0]? arr[409] : arr[408];
wire r1_206;
assign r1_206 = in[0]? arr[411] : arr[410];
wire r1_207;
assign r1_207 = in[0]? arr[413] : arr[412];
wire r1_208;
assign r1_208 = in[0]? arr[415] : arr[414];
wire r1_209;
assign r1_209 = in[0]? arr[417] : arr[416];
wire r1_210;
assign r1_210 = in[0]? arr[419] : arr[418];
wire r1_211;
assign r1_211 = in[0]? arr[421] : arr[420];
wire r1_212;
assign r1_212 = in[0]? arr[423] : arr[422];
wire r1_213;
assign r1_213 = in[0]? arr[425] : arr[424];
wire r1_214;
assign r1_214 = in[0]? arr[427] : arr[426];
wire r1_215;
assign r1_215 = in[0]? arr[429] : arr[428];
wire r1_216;
assign r1_216 = in[0]? arr[431] : arr[430];
wire r1_217;
assign r1_217 = in[0]? arr[433] : arr[432];
wire r1_218;
assign r1_218 = in[0]? arr[435] : arr[434];
wire r1_219;
assign r1_219 = in[0]? arr[437] : arr[436];
wire r1_220;
assign r1_220 = in[0]? arr[439] : arr[438];
wire r1_221;
assign r1_221 = in[0]? arr[441] : arr[440];
wire r1_222;
assign r1_222 = in[0]? arr[443] : arr[442];
wire r1_223;
assign r1_223 = in[0]? arr[445] : arr[444];
wire r1_224;
assign r1_224 = in[0]? arr[447] : arr[446];
wire r1_225;
assign r1_225 = in[0]? arr[449] : arr[448];
wire r1_226;
assign r1_226 = in[0]? arr[451] : arr[450];
wire r1_227;
assign r1_227 = in[0]? arr[453] : arr[452];
wire r1_228;
assign r1_228 = in[0]? arr[455] : arr[454];
wire r1_229;
assign r1_229 = in[0]? arr[457] : arr[456];
wire r1_230;
assign r1_230 = in[0]? arr[459] : arr[458];
wire r1_231;
assign r1_231 = in[0]? arr[461] : arr[460];
wire r1_232;
assign r1_232 = in[0]? arr[463] : arr[462];
wire r1_233;
assign r1_233 = in[0]? arr[465] : arr[464];
wire r1_234;
assign r1_234 = in[0]? arr[467] : arr[466];
wire r1_235;
assign r1_235 = in[0]? arr[469] : arr[468];
wire r1_236;
assign r1_236 = in[0]? arr[471] : arr[470];
wire r1_237;
assign r1_237 = in[0]? arr[473] : arr[472];
wire r1_238;
assign r1_238 = in[0]? arr[475] : arr[474];
wire r1_239;
assign r1_239 = in[0]? arr[477] : arr[476];
wire r1_240;
assign r1_240 = in[0]? arr[479] : arr[478];
wire r1_241;
assign r1_241 = in[0]? arr[481] : arr[480];
wire r1_242;
assign r1_242 = in[0]? arr[483] : arr[482];
wire r1_243;
assign r1_243 = in[0]? arr[485] : arr[484];
wire r1_244;
assign r1_244 = in[0]? arr[487] : arr[486];
wire r1_245;
assign r1_245 = in[0]? arr[489] : arr[488];
wire r1_246;
assign r1_246 = in[0]? arr[491] : arr[490];
wire r1_247;
assign r1_247 = in[0]? arr[493] : arr[492];
wire r1_248;
assign r1_248 = in[0]? arr[495] : arr[494];
wire r1_249;
assign r1_249 = in[0]? arr[497] : arr[496];
wire r1_250;
assign r1_250 = in[0]? arr[499] : arr[498];
wire r1_251;
assign r1_251 = in[0]? arr[501] : arr[500];
wire r1_252;
assign r1_252 = in[0]? arr[503] : arr[502];
wire r1_253;
assign r1_253 = in[0]? arr[505] : arr[504];
wire r1_254;
assign r1_254 = in[0]? arr[507] : arr[506];
wire r1_255;
assign r1_255 = in[0]? arr[509] : arr[508];
wire r1_256;
assign r1_256 = in[0]? arr[511] : arr[510];
wire r1_257;
assign r1_257 = in[0]? arr[513] : arr[512];
wire r1_258;
assign r1_258 = in[0]? arr[515] : arr[514];
wire r1_259;
assign r1_259 = in[0]? arr[517] : arr[516];
wire r1_260;
assign r1_260 = in[0]? arr[519] : arr[518];
wire r1_261;
assign r1_261 = in[0]? arr[521] : arr[520];
wire r1_262;
assign r1_262 = in[0]? arr[523] : arr[522];
wire r1_263;
assign r1_263 = in[0]? arr[525] : arr[524];
wire r1_264;
assign r1_264 = in[0]? arr[527] : arr[526];
wire r1_265;
assign r1_265 = in[0]? arr[529] : arr[528];
wire r1_266;
assign r1_266 = in[0]? arr[531] : arr[530];
wire r1_267;
assign r1_267 = in[0]? arr[533] : arr[532];
wire r1_268;
assign r1_268 = in[0]? arr[535] : arr[534];
wire r1_269;
assign r1_269 = in[0]? arr[537] : arr[536];
wire r1_270;
assign r1_270 = in[0]? arr[539] : arr[538];
wire r1_271;
assign r1_271 = in[0]? arr[541] : arr[540];
wire r1_272;
assign r1_272 = in[0]? arr[543] : arr[542];
wire r1_273;
assign r1_273 = in[0]? arr[545] : arr[544];
wire r1_274;
assign r1_274 = in[0]? arr[547] : arr[546];
wire r1_275;
assign r1_275 = in[0]? arr[549] : arr[548];
wire r1_276;
assign r1_276 = in[0]? arr[551] : arr[550];
wire r1_277;
assign r1_277 = in[0]? arr[553] : arr[552];
wire r1_278;
assign r1_278 = in[0]? arr[555] : arr[554];
wire r1_279;
assign r1_279 = in[0]? arr[557] : arr[556];
wire r1_280;
assign r1_280 = in[0]? arr[559] : arr[558];
wire r1_281;
assign r1_281 = in[0]? arr[561] : arr[560];
wire r1_282;
assign r1_282 = in[0]? arr[563] : arr[562];
wire r1_283;
assign r1_283 = in[0]? arr[565] : arr[564];
wire r1_284;
assign r1_284 = in[0]? arr[567] : arr[566];
wire r1_285;
assign r1_285 = in[0]? arr[569] : arr[568];
wire r1_286;
assign r1_286 = in[0]? arr[571] : arr[570];
wire r1_287;
assign r1_287 = in[0]? arr[573] : arr[572];
wire r1_288;
assign r1_288 = in[0]? arr[575] : arr[574];
wire r1_289;
assign r1_289 = in[0]? arr[577] : arr[576];
wire r1_290;
assign r1_290 = in[0]? arr[579] : arr[578];
wire r1_291;
assign r1_291 = in[0]? arr[581] : arr[580];
wire r1_292;
assign r1_292 = in[0]? arr[583] : arr[582];
wire r1_293;
assign r1_293 = in[0]? arr[585] : arr[584];
wire r1_294;
assign r1_294 = in[0]? arr[587] : arr[586];
wire r1_295;
assign r1_295 = in[0]? arr[589] : arr[588];
wire r1_296;
assign r1_296 = in[0]? arr[591] : arr[590];
wire r1_297;
assign r1_297 = in[0]? arr[593] : arr[592];
wire r1_298;
assign r1_298 = in[0]? arr[595] : arr[594];
wire r1_299;
assign r1_299 = in[0]? arr[597] : arr[596];
wire r1_300;
assign r1_300 = in[0]? arr[599] : arr[598];
wire r1_301;
assign r1_301 = in[0]? arr[601] : arr[600];
wire r1_302;
assign r1_302 = in[0]? arr[603] : arr[602];
wire r1_303;
assign r1_303 = in[0]? arr[605] : arr[604];
wire r1_304;
assign r1_304 = in[0]? arr[607] : arr[606];
wire r1_305;
assign r1_305 = in[0]? arr[609] : arr[608];
wire r1_306;
assign r1_306 = in[0]? arr[611] : arr[610];
wire r1_307;
assign r1_307 = in[0]? arr[613] : arr[612];
wire r1_308;
assign r1_308 = in[0]? arr[615] : arr[614];
wire r1_309;
assign r1_309 = in[0]? arr[617] : arr[616];
wire r1_310;
assign r1_310 = in[0]? arr[619] : arr[618];
wire r1_311;
assign r1_311 = in[0]? arr[621] : arr[620];
wire r1_312;
assign r1_312 = in[0]? arr[623] : arr[622];
wire r1_313;
assign r1_313 = in[0]? arr[625] : arr[624];
wire r1_314;
assign r1_314 = in[0]? arr[627] : arr[626];
wire r1_315;
assign r1_315 = in[0]? arr[629] : arr[628];
wire r1_316;
assign r1_316 = in[0]? arr[631] : arr[630];
wire r1_317;
assign r1_317 = in[0]? arr[633] : arr[632];
wire r1_318;
assign r1_318 = in[0]? arr[635] : arr[634];
wire r1_319;
assign r1_319 = in[0]? arr[637] : arr[636];
wire r1_320;
assign r1_320 = in[0]? arr[639] : arr[638];
wire r1_321;
assign r1_321 = in[0]? arr[641] : arr[640];
wire r1_322;
assign r1_322 = in[0]? arr[643] : arr[642];
wire r1_323;
assign r1_323 = in[0]? arr[645] : arr[644];
wire r1_324;
assign r1_324 = in[0]? arr[647] : arr[646];
wire r1_325;
assign r1_325 = in[0]? arr[649] : arr[648];
wire r1_326;
assign r1_326 = in[0]? arr[651] : arr[650];
wire r1_327;
assign r1_327 = in[0]? arr[653] : arr[652];
wire r1_328;
assign r1_328 = in[0]? arr[655] : arr[654];
wire r1_329;
assign r1_329 = in[0]? arr[657] : arr[656];
wire r1_330;
assign r1_330 = in[0]? arr[659] : arr[658];
wire r1_331;
assign r1_331 = in[0]? arr[661] : arr[660];
wire r1_332;
assign r1_332 = in[0]? arr[663] : arr[662];
wire r1_333;
assign r1_333 = in[0]? arr[665] : arr[664];
wire r1_334;
assign r1_334 = in[0]? arr[667] : arr[666];
wire r1_335;
assign r1_335 = in[0]? arr[669] : arr[668];
wire r1_336;
assign r1_336 = in[0]? arr[671] : arr[670];
wire r1_337;
assign r1_337 = in[0]? arr[673] : arr[672];
wire r1_338;
assign r1_338 = in[0]? arr[675] : arr[674];
wire r1_339;
assign r1_339 = in[0]? arr[677] : arr[676];
wire r1_340;
assign r1_340 = in[0]? arr[679] : arr[678];
wire r1_341;
assign r1_341 = in[0]? arr[681] : arr[680];
wire r1_342;
assign r1_342 = in[0]? arr[683] : arr[682];
wire r1_343;
assign r1_343 = in[0]? arr[685] : arr[684];
wire r1_344;
assign r1_344 = in[0]? arr[687] : arr[686];
wire r1_345;
assign r1_345 = in[0]? arr[689] : arr[688];
wire r1_346;
assign r1_346 = in[0]? arr[691] : arr[690];
wire r1_347;
assign r1_347 = in[0]? arr[693] : arr[692];
wire r1_348;
assign r1_348 = in[0]? arr[695] : arr[694];
wire r1_349;
assign r1_349 = in[0]? arr[697] : arr[696];
wire r1_350;
assign r1_350 = in[0]? arr[699] : arr[698];
wire r1_351;
assign r1_351 = in[0]? arr[701] : arr[700];
wire r1_352;
assign r1_352 = in[0]? arr[703] : arr[702];
wire r1_353;
assign r1_353 = in[0]? arr[705] : arr[704];
wire r1_354;
assign r1_354 = in[0]? arr[707] : arr[706];
wire r1_355;
assign r1_355 = in[0]? arr[709] : arr[708];
wire r1_356;
assign r1_356 = in[0]? arr[711] : arr[710];
wire r1_357;
assign r1_357 = in[0]? arr[713] : arr[712];
wire r1_358;
assign r1_358 = in[0]? arr[715] : arr[714];
wire r1_359;
assign r1_359 = in[0]? arr[717] : arr[716];
wire r1_360;
assign r1_360 = in[0]? arr[719] : arr[718];
wire r1_361;
assign r1_361 = in[0]? arr[721] : arr[720];
wire r1_362;
assign r1_362 = in[0]? arr[723] : arr[722];
wire r1_363;
assign r1_363 = in[0]? arr[725] : arr[724];
wire r1_364;
assign r1_364 = in[0]? arr[727] : arr[726];
wire r1_365;
assign r1_365 = in[0]? arr[729] : arr[728];
wire r1_366;
assign r1_366 = in[0]? arr[731] : arr[730];
wire r1_367;
assign r1_367 = in[0]? arr[733] : arr[732];
wire r1_368;
assign r1_368 = in[0]? arr[735] : arr[734];
wire r1_369;
assign r1_369 = in[0]? arr[737] : arr[736];
wire r1_370;
assign r1_370 = in[0]? arr[739] : arr[738];
wire r1_371;
assign r1_371 = in[0]? arr[741] : arr[740];
wire r1_372;
assign r1_372 = in[0]? arr[743] : arr[742];
wire r1_373;
assign r1_373 = in[0]? arr[745] : arr[744];
wire r1_374;
assign r1_374 = in[0]? arr[747] : arr[746];
wire r1_375;
assign r1_375 = in[0]? arr[749] : arr[748];
wire r1_376;
assign r1_376 = in[0]? arr[751] : arr[750];
wire r1_377;
assign r1_377 = in[0]? arr[753] : arr[752];
wire r1_378;
assign r1_378 = in[0]? arr[755] : arr[754];
wire r1_379;
assign r1_379 = in[0]? arr[757] : arr[756];
wire r1_380;
assign r1_380 = in[0]? arr[759] : arr[758];
wire r1_381;
assign r1_381 = in[0]? arr[761] : arr[760];
wire r1_382;
assign r1_382 = in[0]? arr[763] : arr[762];
wire r1_383;
assign r1_383 = in[0]? arr[765] : arr[764];
wire r1_384;
assign r1_384 = in[0]? arr[767] : arr[766];
wire r1_385;
assign r1_385 = in[0]? arr[769] : arr[768];
wire r1_386;
assign r1_386 = in[0]? arr[771] : arr[770];
wire r1_387;
assign r1_387 = in[0]? arr[773] : arr[772];
wire r1_388;
assign r1_388 = in[0]? arr[775] : arr[774];
wire r1_389;
assign r1_389 = in[0]? arr[777] : arr[776];
wire r1_390;
assign r1_390 = in[0]? arr[779] : arr[778];
wire r1_391;
assign r1_391 = in[0]? arr[781] : arr[780];
wire r1_392;
assign r1_392 = in[0]? arr[783] : arr[782];
wire r1_393;
assign r1_393 = in[0]? arr[785] : arr[784];
wire r1_394;
assign r1_394 = in[0]? arr[787] : arr[786];
wire r1_395;
assign r1_395 = in[0]? arr[789] : arr[788];
wire r1_396;
assign r1_396 = in[0]? arr[791] : arr[790];
wire r1_397;
assign r1_397 = in[0]? arr[793] : arr[792];
wire r1_398;
assign r1_398 = in[0]? arr[795] : arr[794];
wire r1_399;
assign r1_399 = in[0]? arr[797] : arr[796];
wire r1_400;
assign r1_400 = in[0]? arr[799] : arr[798];
wire r1_401;
assign r1_401 = in[0]? arr[801] : arr[800];
wire r1_402;
assign r1_402 = in[0]? arr[803] : arr[802];
wire r1_403;
assign r1_403 = in[0]? arr[805] : arr[804];
wire r1_404;
assign r1_404 = in[0]? arr[807] : arr[806];
wire r1_405;
assign r1_405 = in[0]? arr[809] : arr[808];
wire r1_406;
assign r1_406 = in[0]? arr[811] : arr[810];
wire r1_407;
assign r1_407 = in[0]? arr[813] : arr[812];
wire r1_408;
assign r1_408 = in[0]? arr[815] : arr[814];
wire r1_409;
assign r1_409 = in[0]? arr[817] : arr[816];
wire r1_410;
assign r1_410 = in[0]? arr[819] : arr[818];
wire r1_411;
assign r1_411 = in[0]? arr[821] : arr[820];
wire r1_412;
assign r1_412 = in[0]? arr[823] : arr[822];
wire r1_413;
assign r1_413 = in[0]? arr[825] : arr[824];
wire r1_414;
assign r1_414 = in[0]? arr[827] : arr[826];
wire r1_415;
assign r1_415 = in[0]? arr[829] : arr[828];
wire r1_416;
assign r1_416 = in[0]? arr[831] : arr[830];
wire r1_417;
assign r1_417 = in[0]? arr[833] : arr[832];
wire r1_418;
assign r1_418 = in[0]? arr[835] : arr[834];
wire r1_419;
assign r1_419 = in[0]? arr[837] : arr[836];
wire r1_420;
assign r1_420 = in[0]? arr[839] : arr[838];
wire r1_421;
assign r1_421 = in[0]? arr[841] : arr[840];
wire r1_422;
assign r1_422 = in[0]? arr[843] : arr[842];
wire r1_423;
assign r1_423 = in[0]? arr[845] : arr[844];
wire r1_424;
assign r1_424 = in[0]? arr[847] : arr[846];
wire r1_425;
assign r1_425 = in[0]? arr[849] : arr[848];
wire r1_426;
assign r1_426 = in[0]? arr[851] : arr[850];
wire r1_427;
assign r1_427 = in[0]? arr[853] : arr[852];
wire r1_428;
assign r1_428 = in[0]? arr[855] : arr[854];
wire r1_429;
assign r1_429 = in[0]? arr[857] : arr[856];
wire r1_430;
assign r1_430 = in[0]? arr[859] : arr[858];
wire r1_431;
assign r1_431 = in[0]? arr[861] : arr[860];
wire r1_432;
assign r1_432 = in[0]? arr[863] : arr[862];
wire r1_433;
assign r1_433 = in[0]? arr[865] : arr[864];
wire r1_434;
assign r1_434 = in[0]? arr[867] : arr[866];
wire r1_435;
assign r1_435 = in[0]? arr[869] : arr[868];
wire r1_436;
assign r1_436 = in[0]? arr[871] : arr[870];
wire r1_437;
assign r1_437 = in[0]? arr[873] : arr[872];
wire r1_438;
assign r1_438 = in[0]? arr[875] : arr[874];
wire r1_439;
assign r1_439 = in[0]? arr[877] : arr[876];
wire r1_440;
assign r1_440 = in[0]? arr[879] : arr[878];
wire r1_441;
assign r1_441 = in[0]? arr[881] : arr[880];
wire r1_442;
assign r1_442 = in[0]? arr[883] : arr[882];
wire r1_443;
assign r1_443 = in[0]? arr[885] : arr[884];
wire r1_444;
assign r1_444 = in[0]? arr[887] : arr[886];
wire r1_445;
assign r1_445 = in[0]? arr[889] : arr[888];
wire r1_446;
assign r1_446 = in[0]? arr[891] : arr[890];
wire r1_447;
assign r1_447 = in[0]? arr[893] : arr[892];
wire r1_448;
assign r1_448 = in[0]? arr[895] : arr[894];
wire r1_449;
assign r1_449 = in[0]? arr[897] : arr[896];
wire r1_450;
assign r1_450 = in[0]? arr[899] : arr[898];
wire r1_451;
assign r1_451 = in[0]? arr[901] : arr[900];
wire r1_452;
assign r1_452 = in[0]? arr[903] : arr[902];
wire r1_453;
assign r1_453 = in[0]? arr[905] : arr[904];
wire r1_454;
assign r1_454 = in[0]? arr[907] : arr[906];
wire r1_455;
assign r1_455 = in[0]? arr[909] : arr[908];
wire r1_456;
assign r1_456 = in[0]? arr[911] : arr[910];
wire r1_457;
assign r1_457 = in[0]? arr[913] : arr[912];
wire r1_458;
assign r1_458 = in[0]? arr[915] : arr[914];
wire r1_459;
assign r1_459 = in[0]? arr[917] : arr[916];
wire r1_460;
assign r1_460 = in[0]? arr[919] : arr[918];
wire r1_461;
assign r1_461 = in[0]? arr[921] : arr[920];
wire r1_462;
assign r1_462 = in[0]? arr[923] : arr[922];
wire r1_463;
assign r1_463 = in[0]? arr[925] : arr[924];
wire r1_464;
assign r1_464 = in[0]? arr[927] : arr[926];
wire r1_465;
assign r1_465 = in[0]? arr[929] : arr[928];
wire r1_466;
assign r1_466 = in[0]? arr[931] : arr[930];
wire r1_467;
assign r1_467 = in[0]? arr[933] : arr[932];
wire r1_468;
assign r1_468 = in[0]? arr[935] : arr[934];
wire r1_469;
assign r1_469 = in[0]? arr[937] : arr[936];
wire r1_470;
assign r1_470 = in[0]? arr[939] : arr[938];
wire r1_471;
assign r1_471 = in[0]? arr[941] : arr[940];
wire r1_472;
assign r1_472 = in[0]? arr[943] : arr[942];
wire r1_473;
assign r1_473 = in[0]? arr[945] : arr[944];
wire r1_474;
assign r1_474 = in[0]? arr[947] : arr[946];
wire r1_475;
assign r1_475 = in[0]? arr[949] : arr[948];
wire r1_476;
assign r1_476 = in[0]? arr[951] : arr[950];
wire r1_477;
assign r1_477 = in[0]? arr[953] : arr[952];
wire r1_478;
assign r1_478 = in[0]? arr[955] : arr[954];
wire r1_479;
assign r1_479 = in[0]? arr[957] : arr[956];
wire r1_480;
assign r1_480 = in[0]? arr[959] : arr[958];
wire r1_481;
assign r1_481 = in[0]? arr[961] : arr[960];
wire r1_482;
assign r1_482 = in[0]? arr[963] : arr[962];
wire r1_483;
assign r1_483 = in[0]? arr[965] : arr[964];
wire r1_484;
assign r1_484 = in[0]? arr[967] : arr[966];
wire r1_485;
assign r1_485 = in[0]? arr[969] : arr[968];
wire r1_486;
assign r1_486 = in[0]? arr[971] : arr[970];
wire r1_487;
assign r1_487 = in[0]? arr[973] : arr[972];
wire r1_488;
assign r1_488 = in[0]? arr[975] : arr[974];
wire r1_489;
assign r1_489 = in[0]? arr[977] : arr[976];
wire r1_490;
assign r1_490 = in[0]? arr[979] : arr[978];
wire r1_491;
assign r1_491 = in[0]? arr[981] : arr[980];
wire r1_492;
assign r1_492 = in[0]? arr[983] : arr[982];
wire r1_493;
assign r1_493 = in[0]? arr[985] : arr[984];
wire r1_494;
assign r1_494 = in[0]? arr[987] : arr[986];
wire r1_495;
assign r1_495 = in[0]? arr[989] : arr[988];
wire r1_496;
assign r1_496 = in[0]? arr[991] : arr[990];
wire r1_497;
assign r1_497 = in[0]? arr[993] : arr[992];
wire r1_498;
assign r1_498 = in[0]? arr[995] : arr[994];
wire r1_499;
assign r1_499 = in[0]? arr[997] : arr[996];
wire r1_500;
assign r1_500 = in[0]? arr[999] : arr[998];
wire r1_501;
assign r1_501 = in[0]? arr[1001] : arr[1000];
wire r1_502;
assign r1_502 = in[0]? arr[1003] : arr[1002];
wire r1_503;
assign r1_503 = in[0]? arr[1005] : arr[1004];
wire r1_504;
assign r1_504 = in[0]? arr[1007] : arr[1006];
wire r1_505;
assign r1_505 = in[0]? arr[1009] : arr[1008];
wire r1_506;
assign r1_506 = in[0]? arr[1011] : arr[1010];
wire r1_507;
assign r1_507 = in[0]? arr[1013] : arr[1012];
wire r1_508;
assign r1_508 = in[0]? arr[1015] : arr[1014];
wire r1_509;
assign r1_509 = in[0]? arr[1017] : arr[1016];
wire r1_510;
assign r1_510 = in[0]? arr[1019] : arr[1018];
wire r1_511;
assign r1_511 = in[0]? arr[1021] : arr[1020];
wire r1_512;
assign r1_512 = in[0]? arr[1023] : arr[1022];
wire r1_513;
assign r1_513 = in[0]? arr[1025] : arr[1024];
wire r1_514;
assign r1_514 = in[0]? arr[1027] : arr[1026];
wire r1_515;
assign r1_515 = in[0]? arr[1029] : arr[1028];
wire r1_516;
assign r1_516 = in[0]? arr[1031] : arr[1030];
wire r1_517;
assign r1_517 = in[0]? arr[1033] : arr[1032];
wire r1_518;
assign r1_518 = in[0]? arr[1035] : arr[1034];
wire r1_519;
assign r1_519 = in[0]? arr[1037] : arr[1036];
wire r1_520;
assign r1_520 = in[0]? arr[1039] : arr[1038];
wire r1_521;
assign r1_521 = in[0]? arr[1041] : arr[1040];
wire r1_522;
assign r1_522 = in[0]? arr[1043] : arr[1042];
wire r1_523;
assign r1_523 = in[0]? arr[1045] : arr[1044];
wire r1_524;
assign r1_524 = in[0]? arr[1047] : arr[1046];
wire r1_525;
assign r1_525 = in[0]? arr[1049] : arr[1048];
wire r1_526;
assign r1_526 = in[0]? arr[1051] : arr[1050];
wire r1_527;
assign r1_527 = in[0]? arr[1053] : arr[1052];
wire r1_528;
assign r1_528 = in[0]? arr[1055] : arr[1054];
wire r1_529;
assign r1_529 = in[0]? arr[1057] : arr[1056];
wire r1_530;
assign r1_530 = in[0]? arr[1059] : arr[1058];
wire r1_531;
assign r1_531 = in[0]? arr[1061] : arr[1060];
wire r1_532;
assign r1_532 = in[0]? arr[1063] : arr[1062];
wire r1_533;
assign r1_533 = in[0]? arr[1065] : arr[1064];
wire r1_534;
assign r1_534 = in[0]? arr[1067] : arr[1066];
wire r1_535;
assign r1_535 = in[0]? arr[1069] : arr[1068];
wire r1_536;
assign r1_536 = in[0]? arr[1071] : arr[1070];
wire r1_537;
assign r1_537 = in[0]? arr[1073] : arr[1072];
wire r1_538;
assign r1_538 = in[0]? arr[1075] : arr[1074];
wire r1_539;
assign r1_539 = in[0]? arr[1077] : arr[1076];
wire r1_540;
assign r1_540 = in[0]? arr[1079] : arr[1078];
wire r1_541;
assign r1_541 = in[0]? arr[1081] : arr[1080];
wire r1_542;
assign r1_542 = in[0]? arr[1083] : arr[1082];
wire r1_543;
assign r1_543 = in[0]? arr[1085] : arr[1084];
wire r1_544;
assign r1_544 = in[0]? arr[1087] : arr[1086];
wire r1_545;
assign r1_545 = in[0]? arr[1089] : arr[1088];
wire r1_546;
assign r1_546 = in[0]? arr[1091] : arr[1090];
wire r1_547;
assign r1_547 = in[0]? arr[1093] : arr[1092];
wire r1_548;
assign r1_548 = in[0]? arr[1095] : arr[1094];
wire r1_549;
assign r1_549 = in[0]? arr[1097] : arr[1096];
wire r1_550;
assign r1_550 = in[0]? arr[1099] : arr[1098];
wire r1_551;
assign r1_551 = in[0]? arr[1101] : arr[1100];
wire r1_552;
assign r1_552 = in[0]? arr[1103] : arr[1102];
wire r1_553;
assign r1_553 = in[0]? arr[1105] : arr[1104];
wire r1_554;
assign r1_554 = in[0]? arr[1107] : arr[1106];
wire r1_555;
assign r1_555 = in[0]? arr[1109] : arr[1108];
wire r1_556;
assign r1_556 = in[0]? arr[1111] : arr[1110];
wire r1_557;
assign r1_557 = in[0]? arr[1113] : arr[1112];
wire r1_558;
assign r1_558 = in[0]? arr[1115] : arr[1114];
wire r1_559;
assign r1_559 = in[0]? arr[1117] : arr[1116];
wire r1_560;
assign r1_560 = in[0]? arr[1119] : arr[1118];
wire r1_561;
assign r1_561 = in[0]? arr[1121] : arr[1120];
wire r1_562;
assign r1_562 = in[0]? arr[1123] : arr[1122];
wire r1_563;
assign r1_563 = in[0]? arr[1125] : arr[1124];
wire r1_564;
assign r1_564 = in[0]? arr[1127] : arr[1126];
wire r1_565;
assign r1_565 = in[0]? arr[1129] : arr[1128];
wire r1_566;
assign r1_566 = in[0]? arr[1131] : arr[1130];
wire r1_567;
assign r1_567 = in[0]? arr[1133] : arr[1132];
wire r1_568;
assign r1_568 = in[0]? arr[1135] : arr[1134];
wire r1_569;
assign r1_569 = in[0]? arr[1137] : arr[1136];
wire r1_570;
assign r1_570 = in[0]? arr[1139] : arr[1138];
wire r1_571;
assign r1_571 = in[0]? arr[1141] : arr[1140];
wire r1_572;
assign r1_572 = in[0]? arr[1143] : arr[1142];
wire r1_573;
assign r1_573 = in[0]? arr[1145] : arr[1144];
wire r1_574;
assign r1_574 = in[0]? arr[1147] : arr[1146];
wire r1_575;
assign r1_575 = in[0]? arr[1149] : arr[1148];
wire r1_576;
assign r1_576 = in[0]? arr[1151] : arr[1150];
wire r1_577;
assign r1_577 = in[0]? arr[1153] : arr[1152];
wire r1_578;
assign r1_578 = in[0]? arr[1155] : arr[1154];
wire r1_579;
assign r1_579 = in[0]? arr[1157] : arr[1156];
wire r1_580;
assign r1_580 = in[0]? arr[1159] : arr[1158];
wire r1_581;
assign r1_581 = in[0]? arr[1161] : arr[1160];
wire r1_582;
assign r1_582 = in[0]? arr[1163] : arr[1162];
wire r1_583;
assign r1_583 = in[0]? arr[1165] : arr[1164];
wire r1_584;
assign r1_584 = in[0]? arr[1167] : arr[1166];
wire r1_585;
assign r1_585 = in[0]? arr[1169] : arr[1168];
wire r1_586;
assign r1_586 = in[0]? arr[1171] : arr[1170];
wire r1_587;
assign r1_587 = in[0]? arr[1173] : arr[1172];
wire r1_588;
assign r1_588 = in[0]? arr[1175] : arr[1174];
wire r1_589;
assign r1_589 = in[0]? arr[1177] : arr[1176];
wire r1_590;
assign r1_590 = in[0]? arr[1179] : arr[1178];
wire r1_591;
assign r1_591 = in[0]? arr[1181] : arr[1180];
wire r1_592;
assign r1_592 = in[0]? arr[1183] : arr[1182];
wire r1_593;
assign r1_593 = in[0]? arr[1185] : arr[1184];
wire r1_594;
assign r1_594 = in[0]? arr[1187] : arr[1186];
wire r1_595;
assign r1_595 = in[0]? arr[1189] : arr[1188];
wire r1_596;
assign r1_596 = in[0]? arr[1191] : arr[1190];
wire r1_597;
assign r1_597 = in[0]? arr[1193] : arr[1192];
wire r1_598;
assign r1_598 = in[0]? arr[1195] : arr[1194];
wire r1_599;
assign r1_599 = in[0]? arr[1197] : arr[1196];
wire r1_600;
assign r1_600 = in[0]? arr[1199] : arr[1198];
wire r1_601;
assign r1_601 = in[0]? arr[1201] : arr[1200];
wire r1_602;
assign r1_602 = in[0]? arr[1203] : arr[1202];
wire r1_603;
assign r1_603 = in[0]? arr[1205] : arr[1204];
wire r1_604;
assign r1_604 = in[0]? arr[1207] : arr[1206];
wire r1_605;
assign r1_605 = in[0]? arr[1209] : arr[1208];
wire r1_606;
assign r1_606 = in[0]? arr[1211] : arr[1210];
wire r1_607;
assign r1_607 = in[0]? arr[1213] : arr[1212];
wire r1_608;
assign r1_608 = in[0]? arr[1215] : arr[1214];
wire r1_609;
assign r1_609 = in[0]? arr[1217] : arr[1216];
wire r1_610;
assign r1_610 = in[0]? arr[1219] : arr[1218];
wire r1_611;
assign r1_611 = in[0]? arr[1221] : arr[1220];
wire r1_612;
assign r1_612 = in[0]? arr[1223] : arr[1222];
wire r1_613;
assign r1_613 = in[0]? arr[1225] : arr[1224];
wire r1_614;
assign r1_614 = in[0]? arr[1227] : arr[1226];
wire r1_615;
assign r1_615 = in[0]? arr[1229] : arr[1228];
wire r1_616;
assign r1_616 = in[0]? arr[1231] : arr[1230];
wire r1_617;
assign r1_617 = in[0]? arr[1233] : arr[1232];
wire r1_618;
assign r1_618 = in[0]? arr[1235] : arr[1234];
wire r1_619;
assign r1_619 = in[0]? arr[1237] : arr[1236];
wire r1_620;
assign r1_620 = in[0]? arr[1239] : arr[1238];
wire r1_621;
assign r1_621 = in[0]? arr[1241] : arr[1240];
wire r1_622;
assign r1_622 = in[0]? arr[1243] : arr[1242];
wire r1_623;
assign r1_623 = in[0]? arr[1245] : arr[1244];
wire r1_624;
assign r1_624 = in[0]? arr[1247] : arr[1246];
wire r1_625;
assign r1_625 = in[0]? arr[1249] : arr[1248];
wire r1_626;
assign r1_626 = in[0]? arr[1251] : arr[1250];
wire r1_627;
assign r1_627 = in[0]? arr[1253] : arr[1252];
wire r1_628;
assign r1_628 = in[0]? arr[1255] : arr[1254];
wire r1_629;
assign r1_629 = in[0]? arr[1257] : arr[1256];
wire r1_630;
assign r1_630 = in[0]? arr[1259] : arr[1258];
wire r1_631;
assign r1_631 = in[0]? arr[1261] : arr[1260];
wire r1_632;
assign r1_632 = in[0]? arr[1263] : arr[1262];
wire r1_633;
assign r1_633 = in[0]? arr[1265] : arr[1264];
wire r1_634;
assign r1_634 = in[0]? arr[1267] : arr[1266];
wire r1_635;
assign r1_635 = in[0]? arr[1269] : arr[1268];
wire r1_636;
assign r1_636 = in[0]? arr[1271] : arr[1270];
wire r1_637;
assign r1_637 = in[0]? arr[1273] : arr[1272];
wire r1_638;
assign r1_638 = in[0]? arr[1275] : arr[1274];
wire r1_639;
assign r1_639 = in[0]? arr[1277] : arr[1276];
wire r1_640;
assign r1_640 = in[0]? arr[1279] : arr[1278];
wire r1_641;
assign r1_641 = in[0]? arr[1281] : arr[1280];
wire r1_642;
assign r1_642 = in[0]? arr[1283] : arr[1282];
wire r1_643;
assign r1_643 = in[0]? arr[1285] : arr[1284];
wire r1_644;
assign r1_644 = in[0]? arr[1287] : arr[1286];
wire r1_645;
assign r1_645 = in[0]? arr[1289] : arr[1288];
wire r1_646;
assign r1_646 = in[0]? arr[1291] : arr[1290];
wire r1_647;
assign r1_647 = in[0]? arr[1293] : arr[1292];
wire r1_648;
assign r1_648 = in[0]? arr[1295] : arr[1294];
wire r1_649;
assign r1_649 = in[0]? arr[1297] : arr[1296];
wire r1_650;
assign r1_650 = in[0]? arr[1299] : arr[1298];
wire r1_651;
assign r1_651 = in[0]? arr[1301] : arr[1300];
wire r1_652;
assign r1_652 = in[0]? arr[1303] : arr[1302];
wire r1_653;
assign r1_653 = in[0]? arr[1305] : arr[1304];
wire r1_654;
assign r1_654 = in[0]? arr[1307] : arr[1306];
wire r1_655;
assign r1_655 = in[0]? arr[1309] : arr[1308];
wire r1_656;
assign r1_656 = in[0]? arr[1311] : arr[1310];
wire r1_657;
assign r1_657 = in[0]? arr[1313] : arr[1312];
wire r1_658;
assign r1_658 = in[0]? arr[1315] : arr[1314];
wire r1_659;
assign r1_659 = in[0]? arr[1317] : arr[1316];
wire r1_660;
assign r1_660 = in[0]? arr[1319] : arr[1318];
wire r1_661;
assign r1_661 = in[0]? arr[1321] : arr[1320];
wire r1_662;
assign r1_662 = in[0]? arr[1323] : arr[1322];
wire r1_663;
assign r1_663 = in[0]? arr[1325] : arr[1324];
wire r1_664;
assign r1_664 = in[0]? arr[1327] : arr[1326];
wire r1_665;
assign r1_665 = in[0]? arr[1329] : arr[1328];
wire r1_666;
assign r1_666 = in[0]? arr[1331] : arr[1330];
wire r1_667;
assign r1_667 = in[0]? arr[1333] : arr[1332];
wire r1_668;
assign r1_668 = in[0]? arr[1335] : arr[1334];
wire r1_669;
assign r1_669 = in[0]? arr[1337] : arr[1336];
wire r1_670;
assign r1_670 = in[0]? arr[1339] : arr[1338];
wire r1_671;
assign r1_671 = in[0]? arr[1341] : arr[1340];
wire r1_672;
assign r1_672 = in[0]? arr[1343] : arr[1342];
wire r1_673;
assign r1_673 = in[0]? arr[1345] : arr[1344];
wire r1_674;
assign r1_674 = in[0]? arr[1347] : arr[1346];
wire r1_675;
assign r1_675 = in[0]? arr[1349] : arr[1348];
wire r1_676;
assign r1_676 = in[0]? arr[1351] : arr[1350];
wire r1_677;
assign r1_677 = in[0]? arr[1353] : arr[1352];
wire r1_678;
assign r1_678 = in[0]? arr[1355] : arr[1354];
wire r1_679;
assign r1_679 = in[0]? arr[1357] : arr[1356];
wire r1_680;
assign r1_680 = in[0]? arr[1359] : arr[1358];
wire r1_681;
assign r1_681 = in[0]? arr[1361] : arr[1360];
wire r1_682;
assign r1_682 = in[0]? arr[1363] : arr[1362];
wire r1_683;
assign r1_683 = in[0]? arr[1365] : arr[1364];
wire r1_684;
assign r1_684 = in[0]? arr[1367] : arr[1366];
wire r1_685;
assign r1_685 = in[0]? arr[1369] : arr[1368];
wire r1_686;
assign r1_686 = in[0]? arr[1371] : arr[1370];
wire r1_687;
assign r1_687 = in[0]? arr[1373] : arr[1372];
wire r1_688;
assign r1_688 = in[0]? arr[1375] : arr[1374];
wire r1_689;
assign r1_689 = in[0]? arr[1377] : arr[1376];
wire r1_690;
assign r1_690 = in[0]? arr[1379] : arr[1378];
wire r1_691;
assign r1_691 = in[0]? arr[1381] : arr[1380];
wire r1_692;
assign r1_692 = in[0]? arr[1383] : arr[1382];
wire r1_693;
assign r1_693 = in[0]? arr[1385] : arr[1384];
wire r1_694;
assign r1_694 = in[0]? arr[1387] : arr[1386];
wire r1_695;
assign r1_695 = in[0]? arr[1389] : arr[1388];
wire r1_696;
assign r1_696 = in[0]? arr[1391] : arr[1390];
wire r1_697;
assign r1_697 = in[0]? arr[1393] : arr[1392];
wire r1_698;
assign r1_698 = in[0]? arr[1395] : arr[1394];
wire r1_699;
assign r1_699 = in[0]? arr[1397] : arr[1396];
wire r1_700;
assign r1_700 = in[0]? arr[1399] : arr[1398];
wire r1_701;
assign r1_701 = in[0]? arr[1401] : arr[1400];
wire r1_702;
assign r1_702 = in[0]? arr[1403] : arr[1402];
wire r1_703;
assign r1_703 = in[0]? arr[1405] : arr[1404];
wire r1_704;
assign r1_704 = in[0]? arr[1407] : arr[1406];
wire r1_705;
assign r1_705 = in[0]? arr[1409] : arr[1408];
wire r1_706;
assign r1_706 = in[0]? arr[1411] : arr[1410];
wire r1_707;
assign r1_707 = in[0]? arr[1413] : arr[1412];
wire r1_708;
assign r1_708 = in[0]? arr[1415] : arr[1414];
wire r1_709;
assign r1_709 = in[0]? arr[1417] : arr[1416];
wire r1_710;
assign r1_710 = in[0]? arr[1419] : arr[1418];
wire r1_711;
assign r1_711 = in[0]? arr[1421] : arr[1420];
wire r1_712;
assign r1_712 = in[0]? arr[1423] : arr[1422];
wire r1_713;
assign r1_713 = in[0]? arr[1425] : arr[1424];
wire r1_714;
assign r1_714 = in[0]? arr[1427] : arr[1426];
wire r1_715;
assign r1_715 = in[0]? arr[1429] : arr[1428];
wire r1_716;
assign r1_716 = in[0]? arr[1431] : arr[1430];
wire r1_717;
assign r1_717 = in[0]? arr[1433] : arr[1432];
wire r1_718;
assign r1_718 = in[0]? arr[1435] : arr[1434];
wire r1_719;
assign r1_719 = in[0]? arr[1437] : arr[1436];
wire r1_720;
assign r1_720 = in[0]? arr[1439] : arr[1438];
wire r1_721;
assign r1_721 = in[0]? arr[1441] : arr[1440];
wire r1_722;
assign r1_722 = in[0]? arr[1443] : arr[1442];
wire r1_723;
assign r1_723 = in[0]? arr[1445] : arr[1444];
wire r1_724;
assign r1_724 = in[0]? arr[1447] : arr[1446];
wire r1_725;
assign r1_725 = in[0]? arr[1449] : arr[1448];
wire r1_726;
assign r1_726 = in[0]? arr[1451] : arr[1450];
wire r1_727;
assign r1_727 = in[0]? arr[1453] : arr[1452];
wire r1_728;
assign r1_728 = in[0]? arr[1455] : arr[1454];
wire r1_729;
assign r1_729 = in[0]? arr[1457] : arr[1456];
wire r1_730;
assign r1_730 = in[0]? arr[1459] : arr[1458];
wire r1_731;
assign r1_731 = in[0]? arr[1461] : arr[1460];
wire r1_732;
assign r1_732 = in[0]? arr[1463] : arr[1462];
wire r1_733;
assign r1_733 = in[0]? arr[1465] : arr[1464];
wire r1_734;
assign r1_734 = in[0]? arr[1467] : arr[1466];
wire r1_735;
assign r1_735 = in[0]? arr[1469] : arr[1468];
wire r1_736;
assign r1_736 = in[0]? arr[1471] : arr[1470];
wire r1_737;
assign r1_737 = in[0]? arr[1473] : arr[1472];
wire r1_738;
assign r1_738 = in[0]? arr[1475] : arr[1474];
wire r1_739;
assign r1_739 = in[0]? arr[1477] : arr[1476];
wire r1_740;
assign r1_740 = in[0]? arr[1479] : arr[1478];
wire r1_741;
assign r1_741 = in[0]? arr[1481] : arr[1480];
wire r1_742;
assign r1_742 = in[0]? arr[1483] : arr[1482];
wire r1_743;
assign r1_743 = in[0]? arr[1485] : arr[1484];
wire r1_744;
assign r1_744 = in[0]? arr[1487] : arr[1486];
wire r1_745;
assign r1_745 = in[0]? arr[1489] : arr[1488];
wire r1_746;
assign r1_746 = in[0]? arr[1491] : arr[1490];
wire r1_747;
assign r1_747 = in[0]? arr[1493] : arr[1492];
wire r1_748;
assign r1_748 = in[0]? arr[1495] : arr[1494];
wire r1_749;
assign r1_749 = in[0]? arr[1497] : arr[1496];
wire r1_750;
assign r1_750 = in[0]? arr[1499] : arr[1498];
wire r1_751;
assign r1_751 = in[0]? arr[1501] : arr[1500];
wire r1_752;
assign r1_752 = in[0]? arr[1503] : arr[1502];
wire r1_753;
assign r1_753 = in[0]? arr[1505] : arr[1504];
wire r1_754;
assign r1_754 = in[0]? arr[1507] : arr[1506];
wire r1_755;
assign r1_755 = in[0]? arr[1509] : arr[1508];
wire r1_756;
assign r1_756 = in[0]? arr[1511] : arr[1510];
wire r1_757;
assign r1_757 = in[0]? arr[1513] : arr[1512];
wire r1_758;
assign r1_758 = in[0]? arr[1515] : arr[1514];
wire r1_759;
assign r1_759 = in[0]? arr[1517] : arr[1516];
wire r1_760;
assign r1_760 = in[0]? arr[1519] : arr[1518];
wire r1_761;
assign r1_761 = in[0]? arr[1521] : arr[1520];
wire r1_762;
assign r1_762 = in[0]? arr[1523] : arr[1522];
wire r1_763;
assign r1_763 = in[0]? arr[1525] : arr[1524];
wire r1_764;
assign r1_764 = in[0]? arr[1527] : arr[1526];
wire r1_765;
assign r1_765 = in[0]? arr[1529] : arr[1528];
wire r1_766;
assign r1_766 = in[0]? arr[1531] : arr[1530];
wire r1_767;
assign r1_767 = in[0]? arr[1533] : arr[1532];
wire r1_768;
assign r1_768 = in[0]? arr[1535] : arr[1534];
wire r1_769;
assign r1_769 = in[0]? arr[1537] : arr[1536];
wire r1_770;
assign r1_770 = in[0]? arr[1539] : arr[1538];
wire r1_771;
assign r1_771 = in[0]? arr[1541] : arr[1540];
wire r1_772;
assign r1_772 = in[0]? arr[1543] : arr[1542];
wire r1_773;
assign r1_773 = in[0]? arr[1545] : arr[1544];
wire r1_774;
assign r1_774 = in[0]? arr[1547] : arr[1546];
wire r1_775;
assign r1_775 = in[0]? arr[1549] : arr[1548];
wire r1_776;
assign r1_776 = in[0]? arr[1551] : arr[1550];
wire r1_777;
assign r1_777 = in[0]? arr[1553] : arr[1552];
wire r1_778;
assign r1_778 = in[0]? arr[1555] : arr[1554];
wire r1_779;
assign r1_779 = in[0]? arr[1557] : arr[1556];
wire r1_780;
assign r1_780 = in[0]? arr[1559] : arr[1558];
wire r1_781;
assign r1_781 = in[0]? arr[1561] : arr[1560];
wire r1_782;
assign r1_782 = in[0]? arr[1563] : arr[1562];
wire r1_783;
assign r1_783 = in[0]? arr[1565] : arr[1564];
wire r1_784;
assign r1_784 = in[0]? arr[1567] : arr[1566];
wire r1_785;
assign r1_785 = in[0]? arr[1569] : arr[1568];
wire r1_786;
assign r1_786 = in[0]? arr[1571] : arr[1570];
wire r1_787;
assign r1_787 = in[0]? arr[1573] : arr[1572];
wire r1_788;
assign r1_788 = in[0]? arr[1575] : arr[1574];
wire r1_789;
assign r1_789 = in[0]? arr[1577] : arr[1576];
wire r1_790;
assign r1_790 = in[0]? arr[1579] : arr[1578];
wire r1_791;
assign r1_791 = in[0]? arr[1581] : arr[1580];
wire r1_792;
assign r1_792 = in[0]? arr[1583] : arr[1582];
wire r1_793;
assign r1_793 = in[0]? arr[1585] : arr[1584];
wire r1_794;
assign r1_794 = in[0]? arr[1587] : arr[1586];
wire r1_795;
assign r1_795 = in[0]? arr[1589] : arr[1588];
wire r1_796;
assign r1_796 = in[0]? arr[1591] : arr[1590];
wire r1_797;
assign r1_797 = in[0]? arr[1593] : arr[1592];
wire r1_798;
assign r1_798 = in[0]? arr[1595] : arr[1594];
wire r1_799;
assign r1_799 = in[0]? arr[1597] : arr[1596];
wire r1_800;
assign r1_800 = in[0]? arr[1599] : arr[1598];
wire r1_801;
assign r1_801 = in[0]? arr[1601] : arr[1600];
wire r1_802;
assign r1_802 = in[0]? arr[1603] : arr[1602];
wire r1_803;
assign r1_803 = in[0]? arr[1605] : arr[1604];
wire r1_804;
assign r1_804 = in[0]? arr[1607] : arr[1606];
wire r1_805;
assign r1_805 = in[0]? arr[1609] : arr[1608];
wire r1_806;
assign r1_806 = in[0]? arr[1611] : arr[1610];
wire r1_807;
assign r1_807 = in[0]? arr[1613] : arr[1612];
wire r1_808;
assign r1_808 = in[0]? arr[1615] : arr[1614];
wire r1_809;
assign r1_809 = in[0]? arr[1617] : arr[1616];
wire r1_810;
assign r1_810 = in[0]? arr[1619] : arr[1618];
wire r1_811;
assign r1_811 = in[0]? arr[1621] : arr[1620];
wire r1_812;
assign r1_812 = in[0]? arr[1623] : arr[1622];
wire r1_813;
assign r1_813 = in[0]? arr[1625] : arr[1624];
wire r1_814;
assign r1_814 = in[0]? arr[1627] : arr[1626];
wire r1_815;
assign r1_815 = in[0]? arr[1629] : arr[1628];
wire r1_816;
assign r1_816 = in[0]? arr[1631] : arr[1630];
wire r1_817;
assign r1_817 = in[0]? arr[1633] : arr[1632];
wire r1_818;
assign r1_818 = in[0]? arr[1635] : arr[1634];
wire r1_819;
assign r1_819 = in[0]? arr[1637] : arr[1636];
wire r1_820;
assign r1_820 = in[0]? arr[1639] : arr[1638];
wire r1_821;
assign r1_821 = in[0]? arr[1641] : arr[1640];
wire r1_822;
assign r1_822 = in[0]? arr[1643] : arr[1642];
wire r1_823;
assign r1_823 = in[0]? arr[1645] : arr[1644];
wire r1_824;
assign r1_824 = in[0]? arr[1647] : arr[1646];
wire r1_825;
assign r1_825 = in[0]? arr[1649] : arr[1648];
wire r1_826;
assign r1_826 = in[0]? arr[1651] : arr[1650];
wire r1_827;
assign r1_827 = in[0]? arr[1653] : arr[1652];
wire r1_828;
assign r1_828 = in[0]? arr[1655] : arr[1654];
wire r1_829;
assign r1_829 = in[0]? arr[1657] : arr[1656];
wire r1_830;
assign r1_830 = in[0]? arr[1659] : arr[1658];
wire r1_831;
assign r1_831 = in[0]? arr[1661] : arr[1660];
wire r1_832;
assign r1_832 = in[0]? arr[1663] : arr[1662];
wire r1_833;
assign r1_833 = in[0]? arr[1665] : arr[1664];
wire r1_834;
assign r1_834 = in[0]? arr[1667] : arr[1666];
wire r1_835;
assign r1_835 = in[0]? arr[1669] : arr[1668];
wire r1_836;
assign r1_836 = in[0]? arr[1671] : arr[1670];
wire r1_837;
assign r1_837 = in[0]? arr[1673] : arr[1672];
wire r1_838;
assign r1_838 = in[0]? arr[1675] : arr[1674];
wire r1_839;
assign r1_839 = in[0]? arr[1677] : arr[1676];
wire r1_840;
assign r1_840 = in[0]? arr[1679] : arr[1678];
wire r1_841;
assign r1_841 = in[0]? arr[1681] : arr[1680];
wire r1_842;
assign r1_842 = in[0]? arr[1683] : arr[1682];
wire r1_843;
assign r1_843 = in[0]? arr[1685] : arr[1684];
wire r1_844;
assign r1_844 = in[0]? arr[1687] : arr[1686];
wire r1_845;
assign r1_845 = in[0]? arr[1689] : arr[1688];
wire r1_846;
assign r1_846 = in[0]? arr[1691] : arr[1690];
wire r1_847;
assign r1_847 = in[0]? arr[1693] : arr[1692];
wire r1_848;
assign r1_848 = in[0]? arr[1695] : arr[1694];
wire r1_849;
assign r1_849 = in[0]? arr[1697] : arr[1696];
wire r1_850;
assign r1_850 = in[0]? arr[1699] : arr[1698];
wire r1_851;
assign r1_851 = in[0]? arr[1701] : arr[1700];
wire r1_852;
assign r1_852 = in[0]? arr[1703] : arr[1702];
wire r1_853;
assign r1_853 = in[0]? arr[1705] : arr[1704];
wire r1_854;
assign r1_854 = in[0]? arr[1707] : arr[1706];
wire r1_855;
assign r1_855 = in[0]? arr[1709] : arr[1708];
wire r1_856;
assign r1_856 = in[0]? arr[1711] : arr[1710];
wire r1_857;
assign r1_857 = in[0]? arr[1713] : arr[1712];
wire r1_858;
assign r1_858 = in[0]? arr[1715] : arr[1714];
wire r1_859;
assign r1_859 = in[0]? arr[1717] : arr[1716];
wire r1_860;
assign r1_860 = in[0]? arr[1719] : arr[1718];
wire r1_861;
assign r1_861 = in[0]? arr[1721] : arr[1720];
wire r1_862;
assign r1_862 = in[0]? arr[1723] : arr[1722];
wire r1_863;
assign r1_863 = in[0]? arr[1725] : arr[1724];
wire r1_864;
assign r1_864 = in[0]? arr[1727] : arr[1726];
wire r1_865;
assign r1_865 = in[0]? arr[1729] : arr[1728];
wire r1_866;
assign r1_866 = in[0]? arr[1731] : arr[1730];
wire r1_867;
assign r1_867 = in[0]? arr[1733] : arr[1732];
wire r1_868;
assign r1_868 = in[0]? arr[1735] : arr[1734];
wire r1_869;
assign r1_869 = in[0]? arr[1737] : arr[1736];
wire r1_870;
assign r1_870 = in[0]? arr[1739] : arr[1738];
wire r1_871;
assign r1_871 = in[0]? arr[1741] : arr[1740];
wire r1_872;
assign r1_872 = in[0]? arr[1743] : arr[1742];
wire r1_873;
assign r1_873 = in[0]? arr[1745] : arr[1744];
wire r1_874;
assign r1_874 = in[0]? arr[1747] : arr[1746];
wire r1_875;
assign r1_875 = in[0]? arr[1749] : arr[1748];
wire r1_876;
assign r1_876 = in[0]? arr[1751] : arr[1750];
wire r1_877;
assign r1_877 = in[0]? arr[1753] : arr[1752];
wire r1_878;
assign r1_878 = in[0]? arr[1755] : arr[1754];
wire r1_879;
assign r1_879 = in[0]? arr[1757] : arr[1756];
wire r1_880;
assign r1_880 = in[0]? arr[1759] : arr[1758];
wire r1_881;
assign r1_881 = in[0]? arr[1761] : arr[1760];
wire r1_882;
assign r1_882 = in[0]? arr[1763] : arr[1762];
wire r1_883;
assign r1_883 = in[0]? arr[1765] : arr[1764];
wire r1_884;
assign r1_884 = in[0]? arr[1767] : arr[1766];
wire r1_885;
assign r1_885 = in[0]? arr[1769] : arr[1768];
wire r1_886;
assign r1_886 = in[0]? arr[1771] : arr[1770];
wire r1_887;
assign r1_887 = in[0]? arr[1773] : arr[1772];
wire r1_888;
assign r1_888 = in[0]? arr[1775] : arr[1774];
wire r1_889;
assign r1_889 = in[0]? arr[1777] : arr[1776];
wire r1_890;
assign r1_890 = in[0]? arr[1779] : arr[1778];
wire r1_891;
assign r1_891 = in[0]? arr[1781] : arr[1780];
wire r1_892;
assign r1_892 = in[0]? arr[1783] : arr[1782];
wire r1_893;
assign r1_893 = in[0]? arr[1785] : arr[1784];
wire r1_894;
assign r1_894 = in[0]? arr[1787] : arr[1786];
wire r1_895;
assign r1_895 = in[0]? arr[1789] : arr[1788];
wire r1_896;
assign r1_896 = in[0]? arr[1791] : arr[1790];
wire r1_897;
assign r1_897 = in[0]? arr[1793] : arr[1792];
wire r1_898;
assign r1_898 = in[0]? arr[1795] : arr[1794];
wire r1_899;
assign r1_899 = in[0]? arr[1797] : arr[1796];
wire r1_900;
assign r1_900 = in[0]? arr[1799] : arr[1798];
wire r1_901;
assign r1_901 = in[0]? arr[1801] : arr[1800];
wire r1_902;
assign r1_902 = in[0]? arr[1803] : arr[1802];
wire r1_903;
assign r1_903 = in[0]? arr[1805] : arr[1804];
wire r1_904;
assign r1_904 = in[0]? arr[1807] : arr[1806];
wire r1_905;
assign r1_905 = in[0]? arr[1809] : arr[1808];
wire r1_906;
assign r1_906 = in[0]? arr[1811] : arr[1810];
wire r1_907;
assign r1_907 = in[0]? arr[1813] : arr[1812];
wire r1_908;
assign r1_908 = in[0]? arr[1815] : arr[1814];
wire r1_909;
assign r1_909 = in[0]? arr[1817] : arr[1816];
wire r1_910;
assign r1_910 = in[0]? arr[1819] : arr[1818];
wire r1_911;
assign r1_911 = in[0]? arr[1821] : arr[1820];
wire r1_912;
assign r1_912 = in[0]? arr[1823] : arr[1822];
wire r1_913;
assign r1_913 = in[0]? arr[1825] : arr[1824];
wire r1_914;
assign r1_914 = in[0]? arr[1827] : arr[1826];
wire r1_915;
assign r1_915 = in[0]? arr[1829] : arr[1828];
wire r1_916;
assign r1_916 = in[0]? arr[1831] : arr[1830];
wire r1_917;
assign r1_917 = in[0]? arr[1833] : arr[1832];
wire r1_918;
assign r1_918 = in[0]? arr[1835] : arr[1834];
wire r1_919;
assign r1_919 = in[0]? arr[1837] : arr[1836];
wire r1_920;
assign r1_920 = in[0]? arr[1839] : arr[1838];
wire r1_921;
assign r1_921 = in[0]? arr[1841] : arr[1840];
wire r1_922;
assign r1_922 = in[0]? arr[1843] : arr[1842];
wire r1_923;
assign r1_923 = in[0]? arr[1845] : arr[1844];
wire r1_924;
assign r1_924 = in[0]? arr[1847] : arr[1846];
wire r1_925;
assign r1_925 = in[0]? arr[1849] : arr[1848];
wire r1_926;
assign r1_926 = in[0]? arr[1851] : arr[1850];
wire r1_927;
assign r1_927 = in[0]? arr[1853] : arr[1852];
wire r1_928;
assign r1_928 = in[0]? arr[1855] : arr[1854];
wire r1_929;
assign r1_929 = in[0]? arr[1857] : arr[1856];
wire r1_930;
assign r1_930 = in[0]? arr[1859] : arr[1858];
wire r1_931;
assign r1_931 = in[0]? arr[1861] : arr[1860];
wire r1_932;
assign r1_932 = in[0]? arr[1863] : arr[1862];
wire r1_933;
assign r1_933 = in[0]? arr[1865] : arr[1864];
wire r1_934;
assign r1_934 = in[0]? arr[1867] : arr[1866];
wire r1_935;
assign r1_935 = in[0]? arr[1869] : arr[1868];
wire r1_936;
assign r1_936 = in[0]? arr[1871] : arr[1870];
wire r1_937;
assign r1_937 = in[0]? arr[1873] : arr[1872];
wire r1_938;
assign r1_938 = in[0]? arr[1875] : arr[1874];
wire r1_939;
assign r1_939 = in[0]? arr[1877] : arr[1876];
wire r1_940;
assign r1_940 = in[0]? arr[1879] : arr[1878];
wire r1_941;
assign r1_941 = in[0]? arr[1881] : arr[1880];
wire r1_942;
assign r1_942 = in[0]? arr[1883] : arr[1882];
wire r1_943;
assign r1_943 = in[0]? arr[1885] : arr[1884];
wire r1_944;
assign r1_944 = in[0]? arr[1887] : arr[1886];
wire r1_945;
assign r1_945 = in[0]? arr[1889] : arr[1888];
wire r1_946;
assign r1_946 = in[0]? arr[1891] : arr[1890];
wire r1_947;
assign r1_947 = in[0]? arr[1893] : arr[1892];
wire r1_948;
assign r1_948 = in[0]? arr[1895] : arr[1894];
wire r1_949;
assign r1_949 = in[0]? arr[1897] : arr[1896];
wire r1_950;
assign r1_950 = in[0]? arr[1899] : arr[1898];
wire r1_951;
assign r1_951 = in[0]? arr[1901] : arr[1900];
wire r1_952;
assign r1_952 = in[0]? arr[1903] : arr[1902];
wire r1_953;
assign r1_953 = in[0]? arr[1905] : arr[1904];
wire r1_954;
assign r1_954 = in[0]? arr[1907] : arr[1906];
wire r1_955;
assign r1_955 = in[0]? arr[1909] : arr[1908];
wire r1_956;
assign r1_956 = in[0]? arr[1911] : arr[1910];
wire r1_957;
assign r1_957 = in[0]? arr[1913] : arr[1912];
wire r1_958;
assign r1_958 = in[0]? arr[1915] : arr[1914];
wire r1_959;
assign r1_959 = in[0]? arr[1917] : arr[1916];
wire r1_960;
assign r1_960 = in[0]? arr[1919] : arr[1918];
wire r1_961;
assign r1_961 = in[0]? arr[1921] : arr[1920];
wire r1_962;
assign r1_962 = in[0]? arr[1923] : arr[1922];
wire r1_963;
assign r1_963 = in[0]? arr[1925] : arr[1924];
wire r1_964;
assign r1_964 = in[0]? arr[1927] : arr[1926];
wire r1_965;
assign r1_965 = in[0]? arr[1929] : arr[1928];
wire r1_966;
assign r1_966 = in[0]? arr[1931] : arr[1930];
wire r1_967;
assign r1_967 = in[0]? arr[1933] : arr[1932];
wire r1_968;
assign r1_968 = in[0]? arr[1935] : arr[1934];
wire r1_969;
assign r1_969 = in[0]? arr[1937] : arr[1936];
wire r1_970;
assign r1_970 = in[0]? arr[1939] : arr[1938];
wire r1_971;
assign r1_971 = in[0]? arr[1941] : arr[1940];
wire r1_972;
assign r1_972 = in[0]? arr[1943] : arr[1942];
wire r1_973;
assign r1_973 = in[0]? arr[1945] : arr[1944];
wire r1_974;
assign r1_974 = in[0]? arr[1947] : arr[1946];
wire r1_975;
assign r1_975 = in[0]? arr[1949] : arr[1948];
wire r1_976;
assign r1_976 = in[0]? arr[1951] : arr[1950];
wire r1_977;
assign r1_977 = in[0]? arr[1953] : arr[1952];
wire r1_978;
assign r1_978 = in[0]? arr[1955] : arr[1954];
wire r1_979;
assign r1_979 = in[0]? arr[1957] : arr[1956];
wire r1_980;
assign r1_980 = in[0]? arr[1959] : arr[1958];
wire r1_981;
assign r1_981 = in[0]? arr[1961] : arr[1960];
wire r1_982;
assign r1_982 = in[0]? arr[1963] : arr[1962];
wire r1_983;
assign r1_983 = in[0]? arr[1965] : arr[1964];
wire r1_984;
assign r1_984 = in[0]? arr[1967] : arr[1966];
wire r1_985;
assign r1_985 = in[0]? arr[1969] : arr[1968];
wire r1_986;
assign r1_986 = in[0]? arr[1971] : arr[1970];
wire r1_987;
assign r1_987 = in[0]? arr[1973] : arr[1972];
wire r1_988;
assign r1_988 = in[0]? arr[1975] : arr[1974];
wire r1_989;
assign r1_989 = in[0]? arr[1977] : arr[1976];
wire r1_990;
assign r1_990 = in[0]? arr[1979] : arr[1978];
wire r1_991;
assign r1_991 = in[0]? arr[1981] : arr[1980];
wire r1_992;
assign r1_992 = in[0]? arr[1983] : arr[1982];
wire r1_993;
assign r1_993 = in[0]? arr[1985] : arr[1984];
wire r1_994;
assign r1_994 = in[0]? arr[1987] : arr[1986];
wire r1_995;
assign r1_995 = in[0]? arr[1989] : arr[1988];
wire r1_996;
assign r1_996 = in[0]? arr[1991] : arr[1990];
wire r1_997;
assign r1_997 = in[0]? arr[1993] : arr[1992];
wire r1_998;
assign r1_998 = in[0]? arr[1995] : arr[1994];
wire r1_999;
assign r1_999 = in[0]? arr[1997] : arr[1996];
wire r1_1000;
assign r1_1000 = in[0]? arr[1999] : arr[1998];
wire r1_1001;
assign r1_1001 = in[0]? arr[2001] : arr[2000];
wire r1_1002;
assign r1_1002 = in[0]? arr[2003] : arr[2002];
wire r1_1003;
assign r1_1003 = in[0]? arr[2005] : arr[2004];
wire r1_1004;
assign r1_1004 = in[0]? arr[2007] : arr[2006];
wire r1_1005;
assign r1_1005 = in[0]? arr[2009] : arr[2008];
wire r1_1006;
assign r1_1006 = in[0]? arr[2011] : arr[2010];
wire r1_1007;
assign r1_1007 = in[0]? arr[2013] : arr[2012];
wire r1_1008;
assign r1_1008 = in[0]? arr[2015] : arr[2014];
wire r1_1009;
assign r1_1009 = in[0]? arr[2017] : arr[2016];
wire r1_1010;
assign r1_1010 = in[0]? arr[2019] : arr[2018];
wire r1_1011;
assign r1_1011 = in[0]? arr[2021] : arr[2020];
wire r1_1012;
assign r1_1012 = in[0]? arr[2023] : arr[2022];
wire r1_1013;
assign r1_1013 = in[0]? arr[2025] : arr[2024];
wire r1_1014;
assign r1_1014 = in[0]? arr[2027] : arr[2026];
wire r1_1015;
assign r1_1015 = in[0]? arr[2029] : arr[2028];
wire r1_1016;
assign r1_1016 = in[0]? arr[2031] : arr[2030];
wire r1_1017;
assign r1_1017 = in[0]? arr[2033] : arr[2032];
wire r1_1018;
assign r1_1018 = in[0]? arr[2035] : arr[2034];
wire r1_1019;
assign r1_1019 = in[0]? arr[2037] : arr[2036];
wire r1_1020;
assign r1_1020 = in[0]? arr[2039] : arr[2038];
wire r1_1021;
assign r1_1021 = in[0]? arr[2041] : arr[2040];
wire r1_1022;
assign r1_1022 = in[0]? arr[2043] : arr[2042];
wire r1_1023;
assign r1_1023 = in[0]? arr[2045] : arr[2044];
wire r1_1024;
assign r1_1024 = in[0]? arr[2047] : arr[2046];
wire r1_1025;
assign r1_1025 = in[0]? arr[2049] : arr[2048];
wire r1_1026;
assign r1_1026 = in[0]? arr[2051] : arr[2050];
wire r1_1027;
assign r1_1027 = in[0]? arr[2053] : arr[2052];
wire r1_1028;
assign r1_1028 = in[0]? arr[2055] : arr[2054];
wire r1_1029;
assign r1_1029 = in[0]? arr[2057] : arr[2056];
wire r1_1030;
assign r1_1030 = in[0]? arr[2059] : arr[2058];
wire r1_1031;
assign r1_1031 = in[0]? arr[2061] : arr[2060];
wire r1_1032;
assign r1_1032 = in[0]? arr[2063] : arr[2062];
wire r1_1033;
assign r1_1033 = in[0]? arr[2065] : arr[2064];
wire r1_1034;
assign r1_1034 = in[0]? arr[2067] : arr[2066];
wire r1_1035;
assign r1_1035 = in[0]? arr[2069] : arr[2068];
wire r1_1036;
assign r1_1036 = in[0]? arr[2071] : arr[2070];
wire r1_1037;
assign r1_1037 = in[0]? arr[2073] : arr[2072];
wire r1_1038;
assign r1_1038 = in[0]? arr[2075] : arr[2074];
wire r1_1039;
assign r1_1039 = in[0]? arr[2077] : arr[2076];
wire r1_1040;
assign r1_1040 = in[0]? arr[2079] : arr[2078];
wire r1_1041;
assign r1_1041 = in[0]? arr[2081] : arr[2080];
wire r1_1042;
assign r1_1042 = in[0]? arr[2083] : arr[2082];
wire r1_1043;
assign r1_1043 = in[0]? arr[2085] : arr[2084];
wire r1_1044;
assign r1_1044 = in[0]? arr[2087] : arr[2086];
wire r1_1045;
assign r1_1045 = in[0]? arr[2089] : arr[2088];
wire r1_1046;
assign r1_1046 = in[0]? arr[2091] : arr[2090];
wire r1_1047;
assign r1_1047 = in[0]? arr[2093] : arr[2092];
wire r1_1048;
assign r1_1048 = in[0]? arr[2095] : arr[2094];
wire r1_1049;
assign r1_1049 = in[0]? arr[2097] : arr[2096];
wire r1_1050;
assign r1_1050 = in[0]? arr[2099] : arr[2098];
wire r1_1051;
assign r1_1051 = in[0]? arr[2101] : arr[2100];
wire r1_1052;
assign r1_1052 = in[0]? arr[2103] : arr[2102];
wire r1_1053;
assign r1_1053 = in[0]? arr[2105] : arr[2104];
wire r1_1054;
assign r1_1054 = in[0]? arr[2107] : arr[2106];
wire r1_1055;
assign r1_1055 = in[0]? arr[2109] : arr[2108];
wire r1_1056;
assign r1_1056 = in[0]? arr[2111] : arr[2110];
wire r1_1057;
assign r1_1057 = in[0]? arr[2113] : arr[2112];
wire r1_1058;
assign r1_1058 = in[0]? arr[2115] : arr[2114];
wire r1_1059;
assign r1_1059 = in[0]? arr[2117] : arr[2116];
wire r1_1060;
assign r1_1060 = in[0]? arr[2119] : arr[2118];
wire r1_1061;
assign r1_1061 = in[0]? arr[2121] : arr[2120];
wire r1_1062;
assign r1_1062 = in[0]? arr[2123] : arr[2122];
wire r1_1063;
assign r1_1063 = in[0]? arr[2125] : arr[2124];
wire r1_1064;
assign r1_1064 = in[0]? arr[2127] : arr[2126];
wire r1_1065;
assign r1_1065 = in[0]? arr[2129] : arr[2128];
wire r1_1066;
assign r1_1066 = in[0]? arr[2131] : arr[2130];
wire r1_1067;
assign r1_1067 = in[0]? arr[2133] : arr[2132];
wire r1_1068;
assign r1_1068 = in[0]? arr[2135] : arr[2134];
wire r1_1069;
assign r1_1069 = in[0]? arr[2137] : arr[2136];
wire r1_1070;
assign r1_1070 = in[0]? arr[2139] : arr[2138];
wire r1_1071;
assign r1_1071 = in[0]? arr[2141] : arr[2140];
wire r1_1072;
assign r1_1072 = in[0]? arr[2143] : arr[2142];
wire r1_1073;
assign r1_1073 = in[0]? arr[2145] : arr[2144];
wire r1_1074;
assign r1_1074 = in[0]? arr[2147] : arr[2146];
wire r1_1075;
assign r1_1075 = in[0]? arr[2149] : arr[2148];
wire r1_1076;
assign r1_1076 = in[0]? arr[2151] : arr[2150];
wire r1_1077;
assign r1_1077 = in[0]? arr[2153] : arr[2152];
wire r1_1078;
assign r1_1078 = in[0]? arr[2155] : arr[2154];
wire r1_1079;
assign r1_1079 = in[0]? arr[2157] : arr[2156];
wire r1_1080;
assign r1_1080 = in[0]? arr[2159] : arr[2158];
wire r1_1081;
assign r1_1081 = in[0]? arr[2161] : arr[2160];
wire r1_1082;
assign r1_1082 = in[0]? arr[2163] : arr[2162];
wire r1_1083;
assign r1_1083 = in[0]? arr[2165] : arr[2164];
wire r1_1084;
assign r1_1084 = in[0]? arr[2167] : arr[2166];
wire r1_1085;
assign r1_1085 = in[0]? arr[2169] : arr[2168];
wire r1_1086;
assign r1_1086 = in[0]? arr[2171] : arr[2170];
wire r1_1087;
assign r1_1087 = in[0]? arr[2173] : arr[2172];
wire r1_1088;
assign r1_1088 = in[0]? arr[2175] : arr[2174];
wire r1_1089;
assign r1_1089 = in[0]? arr[2177] : arr[2176];
wire r1_1090;
assign r1_1090 = in[0]? arr[2179] : arr[2178];
wire r1_1091;
assign r1_1091 = in[0]? arr[2181] : arr[2180];
wire r1_1092;
assign r1_1092 = in[0]? arr[2183] : arr[2182];
wire r1_1093;
assign r1_1093 = in[0]? arr[2185] : arr[2184];
wire r1_1094;
assign r1_1094 = in[0]? arr[2187] : arr[2186];
wire r1_1095;
assign r1_1095 = in[0]? arr[2189] : arr[2188];
wire r1_1096;
assign r1_1096 = in[0]? arr[2191] : arr[2190];
wire r1_1097;
assign r1_1097 = in[0]? arr[2193] : arr[2192];
wire r1_1098;
assign r1_1098 = in[0]? arr[2195] : arr[2194];
wire r1_1099;
assign r1_1099 = in[0]? arr[2197] : arr[2196];
wire r1_1100;
assign r1_1100 = in[0]? arr[2199] : arr[2198];
wire r1_1101;
assign r1_1101 = in[0]? arr[2201] : arr[2200];
wire r1_1102;
assign r1_1102 = in[0]? arr[2203] : arr[2202];
wire r1_1103;
assign r1_1103 = in[0]? arr[2205] : arr[2204];
wire r1_1104;
assign r1_1104 = in[0]? arr[2207] : arr[2206];
wire r1_1105;
assign r1_1105 = in[0]? arr[2209] : arr[2208];
wire r1_1106;
assign r1_1106 = in[0]? arr[2211] : arr[2210];
wire r1_1107;
assign r1_1107 = in[0]? arr[2213] : arr[2212];
wire r1_1108;
assign r1_1108 = in[0]? arr[2215] : arr[2214];
wire r1_1109;
assign r1_1109 = in[0]? arr[2217] : arr[2216];
wire r1_1110;
assign r1_1110 = in[0]? arr[2219] : arr[2218];
wire r1_1111;
assign r1_1111 = in[0]? arr[2221] : arr[2220];
wire r1_1112;
assign r1_1112 = in[0]? arr[2223] : arr[2222];
wire r1_1113;
assign r1_1113 = in[0]? arr[2225] : arr[2224];
wire r1_1114;
assign r1_1114 = in[0]? arr[2227] : arr[2226];
wire r1_1115;
assign r1_1115 = in[0]? arr[2229] : arr[2228];
wire r1_1116;
assign r1_1116 = in[0]? arr[2231] : arr[2230];
wire r1_1117;
assign r1_1117 = in[0]? arr[2233] : arr[2232];
wire r1_1118;
assign r1_1118 = in[0]? arr[2235] : arr[2234];
wire r1_1119;
assign r1_1119 = in[0]? arr[2237] : arr[2236];
wire r1_1120;
assign r1_1120 = in[0]? arr[2239] : arr[2238];
wire r1_1121;
assign r1_1121 = in[0]? arr[2241] : arr[2240];
wire r1_1122;
assign r1_1122 = in[0]? arr[2243] : arr[2242];
wire r1_1123;
assign r1_1123 = in[0]? arr[2245] : arr[2244];
wire r1_1124;
assign r1_1124 = in[0]? arr[2247] : arr[2246];
wire r1_1125;
assign r1_1125 = in[0]? arr[2249] : arr[2248];
wire r1_1126;
assign r1_1126 = in[0]? arr[2251] : arr[2250];
wire r1_1127;
assign r1_1127 = in[0]? arr[2253] : arr[2252];
wire r1_1128;
assign r1_1128 = in[0]? arr[2255] : arr[2254];
wire r1_1129;
assign r1_1129 = in[0]? arr[2257] : arr[2256];
wire r1_1130;
assign r1_1130 = in[0]? arr[2259] : arr[2258];
wire r1_1131;
assign r1_1131 = in[0]? arr[2261] : arr[2260];
wire r1_1132;
assign r1_1132 = in[0]? arr[2263] : arr[2262];
wire r1_1133;
assign r1_1133 = in[0]? arr[2265] : arr[2264];
wire r1_1134;
assign r1_1134 = in[0]? arr[2267] : arr[2266];
wire r1_1135;
assign r1_1135 = in[0]? arr[2269] : arr[2268];
wire r1_1136;
assign r1_1136 = in[0]? arr[2271] : arr[2270];
wire r1_1137;
assign r1_1137 = in[0]? arr[2273] : arr[2272];
wire r1_1138;
assign r1_1138 = in[0]? arr[2275] : arr[2274];
wire r1_1139;
assign r1_1139 = in[0]? arr[2277] : arr[2276];
wire r1_1140;
assign r1_1140 = in[0]? arr[2279] : arr[2278];
wire r1_1141;
assign r1_1141 = in[0]? arr[2281] : arr[2280];
wire r1_1142;
assign r1_1142 = in[0]? arr[2283] : arr[2282];
wire r1_1143;
assign r1_1143 = in[0]? arr[2285] : arr[2284];
wire r1_1144;
assign r1_1144 = in[0]? arr[2287] : arr[2286];
wire r1_1145;
assign r1_1145 = in[0]? arr[2289] : arr[2288];
wire r1_1146;
assign r1_1146 = in[0]? arr[2291] : arr[2290];
wire r1_1147;
assign r1_1147 = in[0]? arr[2293] : arr[2292];
wire r1_1148;
assign r1_1148 = in[0]? arr[2295] : arr[2294];
wire r1_1149;
assign r1_1149 = in[0]? arr[2297] : arr[2296];
wire r1_1150;
assign r1_1150 = in[0]? arr[2299] : arr[2298];
wire r1_1151;
assign r1_1151 = in[0]? arr[2301] : arr[2300];
wire r1_1152;
assign r1_1152 = in[0]? arr[2303] : arr[2302];
wire r1_1153;
assign r1_1153 = in[0]? arr[2305] : arr[2304];
wire r1_1154;
assign r1_1154 = in[0]? arr[2307] : arr[2306];
wire r1_1155;
assign r1_1155 = in[0]? arr[2309] : arr[2308];
wire r1_1156;
assign r1_1156 = in[0]? arr[2311] : arr[2310];
wire r1_1157;
assign r1_1157 = in[0]? arr[2313] : arr[2312];
wire r1_1158;
assign r1_1158 = in[0]? arr[2315] : arr[2314];
wire r1_1159;
assign r1_1159 = in[0]? arr[2317] : arr[2316];
wire r1_1160;
assign r1_1160 = in[0]? arr[2319] : arr[2318];
wire r1_1161;
assign r1_1161 = in[0]? arr[2321] : arr[2320];
wire r1_1162;
assign r1_1162 = in[0]? arr[2323] : arr[2322];
wire r1_1163;
assign r1_1163 = in[0]? arr[2325] : arr[2324];
wire r1_1164;
assign r1_1164 = in[0]? arr[2327] : arr[2326];
wire r1_1165;
assign r1_1165 = in[0]? arr[2329] : arr[2328];
wire r1_1166;
assign r1_1166 = in[0]? arr[2331] : arr[2330];
wire r1_1167;
assign r1_1167 = in[0]? arr[2333] : arr[2332];
wire r1_1168;
assign r1_1168 = in[0]? arr[2335] : arr[2334];
wire r1_1169;
assign r1_1169 = in[0]? arr[2337] : arr[2336];
wire r1_1170;
assign r1_1170 = in[0]? arr[2339] : arr[2338];
wire r1_1171;
assign r1_1171 = in[0]? arr[2341] : arr[2340];
wire r1_1172;
assign r1_1172 = in[0]? arr[2343] : arr[2342];
wire r1_1173;
assign r1_1173 = in[0]? arr[2345] : arr[2344];
wire r1_1174;
assign r1_1174 = in[0]? arr[2347] : arr[2346];
wire r1_1175;
assign r1_1175 = in[0]? arr[2349] : arr[2348];
wire r1_1176;
assign r1_1176 = in[0]? arr[2351] : arr[2350];
wire r1_1177;
assign r1_1177 = in[0]? arr[2353] : arr[2352];
wire r1_1178;
assign r1_1178 = in[0]? arr[2355] : arr[2354];
wire r1_1179;
assign r1_1179 = in[0]? arr[2357] : arr[2356];
wire r1_1180;
assign r1_1180 = in[0]? arr[2359] : arr[2358];
wire r1_1181;
assign r1_1181 = in[0]? arr[2361] : arr[2360];
wire r1_1182;
assign r1_1182 = in[0]? arr[2363] : arr[2362];
wire r1_1183;
assign r1_1183 = in[0]? arr[2365] : arr[2364];
wire r1_1184;
assign r1_1184 = in[0]? arr[2367] : arr[2366];
wire r1_1185;
assign r1_1185 = in[0]? arr[2369] : arr[2368];
wire r1_1186;
assign r1_1186 = in[0]? arr[2371] : arr[2370];
wire r1_1187;
assign r1_1187 = in[0]? arr[2373] : arr[2372];
wire r1_1188;
assign r1_1188 = in[0]? arr[2375] : arr[2374];
wire r1_1189;
assign r1_1189 = in[0]? arr[2377] : arr[2376];
wire r1_1190;
assign r1_1190 = in[0]? arr[2379] : arr[2378];
wire r1_1191;
assign r1_1191 = in[0]? arr[2381] : arr[2380];
wire r1_1192;
assign r1_1192 = in[0]? arr[2383] : arr[2382];
wire r1_1193;
assign r1_1193 = in[0]? arr[2385] : arr[2384];
wire r1_1194;
assign r1_1194 = in[0]? arr[2387] : arr[2386];
wire r1_1195;
assign r1_1195 = in[0]? arr[2389] : arr[2388];
wire r1_1196;
assign r1_1196 = in[0]? arr[2391] : arr[2390];
wire r1_1197;
assign r1_1197 = in[0]? arr[2393] : arr[2392];
wire r1_1198;
assign r1_1198 = in[0]? arr[2395] : arr[2394];
wire r1_1199;
assign r1_1199 = in[0]? arr[2397] : arr[2396];
wire r1_1200;
assign r1_1200 = in[0]? arr[2399] : arr[2398];
wire r1_1201;
assign r1_1201 = in[0]? arr[2401] : arr[2400];
wire r1_1202;
assign r1_1202 = in[0]? arr[2403] : arr[2402];
wire r1_1203;
assign r1_1203 = in[0]? arr[2405] : arr[2404];
wire r1_1204;
assign r1_1204 = in[0]? arr[2407] : arr[2406];
wire r1_1205;
assign r1_1205 = in[0]? arr[2409] : arr[2408];
wire r1_1206;
assign r1_1206 = in[0]? arr[2411] : arr[2410];
wire r1_1207;
assign r1_1207 = in[0]? arr[2413] : arr[2412];
wire r1_1208;
assign r1_1208 = in[0]? arr[2415] : arr[2414];
wire r1_1209;
assign r1_1209 = in[0]? arr[2417] : arr[2416];
wire r1_1210;
assign r1_1210 = in[0]? arr[2419] : arr[2418];
wire r1_1211;
assign r1_1211 = in[0]? arr[2421] : arr[2420];
wire r1_1212;
assign r1_1212 = in[0]? arr[2423] : arr[2422];
wire r1_1213;
assign r1_1213 = in[0]? arr[2425] : arr[2424];
wire r1_1214;
assign r1_1214 = in[0]? arr[2427] : arr[2426];
wire r1_1215;
assign r1_1215 = in[0]? arr[2429] : arr[2428];
wire r1_1216;
assign r1_1216 = in[0]? arr[2431] : arr[2430];
wire r1_1217;
assign r1_1217 = in[0]? arr[2433] : arr[2432];
wire r1_1218;
assign r1_1218 = in[0]? arr[2435] : arr[2434];
wire r1_1219;
assign r1_1219 = in[0]? arr[2437] : arr[2436];
wire r1_1220;
assign r1_1220 = in[0]? arr[2439] : arr[2438];
wire r1_1221;
assign r1_1221 = in[0]? arr[2441] : arr[2440];
wire r1_1222;
assign r1_1222 = in[0]? arr[2443] : arr[2442];
wire r1_1223;
assign r1_1223 = in[0]? arr[2445] : arr[2444];
wire r1_1224;
assign r1_1224 = in[0]? arr[2447] : arr[2446];
wire r1_1225;
assign r1_1225 = in[0]? arr[2449] : arr[2448];
wire r1_1226;
assign r1_1226 = in[0]? arr[2451] : arr[2450];
wire r1_1227;
assign r1_1227 = in[0]? arr[2453] : arr[2452];
wire r1_1228;
assign r1_1228 = in[0]? arr[2455] : arr[2454];
wire r1_1229;
assign r1_1229 = in[0]? arr[2457] : arr[2456];
wire r1_1230;
assign r1_1230 = in[0]? arr[2459] : arr[2458];
wire r1_1231;
assign r1_1231 = in[0]? arr[2461] : arr[2460];
wire r1_1232;
assign r1_1232 = in[0]? arr[2463] : arr[2462];
wire r1_1233;
assign r1_1233 = in[0]? arr[2465] : arr[2464];
wire r1_1234;
assign r1_1234 = in[0]? arr[2467] : arr[2466];
wire r1_1235;
assign r1_1235 = in[0]? arr[2469] : arr[2468];
wire r1_1236;
assign r1_1236 = in[0]? arr[2471] : arr[2470];
wire r1_1237;
assign r1_1237 = in[0]? arr[2473] : arr[2472];
wire r1_1238;
assign r1_1238 = in[0]? arr[2475] : arr[2474];
wire r1_1239;
assign r1_1239 = in[0]? arr[2477] : arr[2476];
wire r1_1240;
assign r1_1240 = in[0]? arr[2479] : arr[2478];
wire r1_1241;
assign r1_1241 = in[0]? arr[2481] : arr[2480];
wire r1_1242;
assign r1_1242 = in[0]? arr[2483] : arr[2482];
wire r1_1243;
assign r1_1243 = in[0]? arr[2485] : arr[2484];
wire r1_1244;
assign r1_1244 = in[0]? arr[2487] : arr[2486];
wire r1_1245;
assign r1_1245 = in[0]? arr[2489] : arr[2488];
wire r1_1246;
assign r1_1246 = in[0]? arr[2491] : arr[2490];
wire r1_1247;
assign r1_1247 = in[0]? arr[2493] : arr[2492];
wire r1_1248;
assign r1_1248 = in[0]? arr[2495] : arr[2494];
wire r1_1249;
assign r1_1249 = in[0]? arr[2497] : arr[2496];
wire r1_1250;
assign r1_1250 = in[0]? arr[2499] : arr[2498];
wire r1_1251;
assign r1_1251 = in[0]? arr[2501] : arr[2500];
wire r1_1252;
assign r1_1252 = in[0]? arr[2503] : arr[2502];
wire r1_1253;
assign r1_1253 = in[0]? arr[2505] : arr[2504];
wire r1_1254;
assign r1_1254 = in[0]? arr[2507] : arr[2506];
wire r1_1255;
assign r1_1255 = in[0]? arr[2509] : arr[2508];
wire r1_1256;
assign r1_1256 = in[0]? arr[2511] : arr[2510];
wire r1_1257;
assign r1_1257 = in[0]? arr[2513] : arr[2512];
wire r1_1258;
assign r1_1258 = in[0]? arr[2515] : arr[2514];
wire r1_1259;
assign r1_1259 = in[0]? arr[2517] : arr[2516];
wire r1_1260;
assign r1_1260 = in[0]? arr[2519] : arr[2518];
wire r1_1261;
assign r1_1261 = in[0]? arr[2521] : arr[2520];
wire r1_1262;
assign r1_1262 = in[0]? arr[2523] : arr[2522];
wire r1_1263;
assign r1_1263 = in[0]? arr[2525] : arr[2524];
wire r1_1264;
assign r1_1264 = in[0]? arr[2527] : arr[2526];
wire r1_1265;
assign r1_1265 = in[0]? arr[2529] : arr[2528];
wire r1_1266;
assign r1_1266 = in[0]? arr[2531] : arr[2530];
wire r1_1267;
assign r1_1267 = in[0]? arr[2533] : arr[2532];
wire r1_1268;
assign r1_1268 = in[0]? arr[2535] : arr[2534];
wire r1_1269;
assign r1_1269 = in[0]? arr[2537] : arr[2536];
wire r1_1270;
assign r1_1270 = in[0]? arr[2539] : arr[2538];
wire r1_1271;
assign r1_1271 = in[0]? arr[2541] : arr[2540];
wire r1_1272;
assign r1_1272 = in[0]? arr[2543] : arr[2542];
wire r1_1273;
assign r1_1273 = in[0]? arr[2545] : arr[2544];
wire r1_1274;
assign r1_1274 = in[0]? arr[2547] : arr[2546];
wire r1_1275;
assign r1_1275 = in[0]? arr[2549] : arr[2548];
wire r1_1276;
assign r1_1276 = in[0]? arr[2551] : arr[2550];
wire r1_1277;
assign r1_1277 = in[0]? arr[2553] : arr[2552];
wire r1_1278;
assign r1_1278 = in[0]? arr[2555] : arr[2554];
wire r1_1279;
assign r1_1279 = in[0]? arr[2557] : arr[2556];
wire r1_1280;
assign r1_1280 = in[0]? arr[2559] : arr[2558];
wire r1_1281;
assign r1_1281 = in[0]? arr[2561] : arr[2560];
wire r1_1282;
assign r1_1282 = in[0]? arr[2563] : arr[2562];
wire r1_1283;
assign r1_1283 = in[0]? arr[2565] : arr[2564];
wire r1_1284;
assign r1_1284 = in[0]? arr[2567] : arr[2566];
wire r1_1285;
assign r1_1285 = in[0]? arr[2569] : arr[2568];
wire r1_1286;
assign r1_1286 = in[0]? arr[2571] : arr[2570];
wire r1_1287;
assign r1_1287 = in[0]? arr[2573] : arr[2572];
wire r1_1288;
assign r1_1288 = in[0]? arr[2575] : arr[2574];
wire r1_1289;
assign r1_1289 = in[0]? arr[2577] : arr[2576];
wire r1_1290;
assign r1_1290 = in[0]? arr[2579] : arr[2578];
wire r1_1291;
assign r1_1291 = in[0]? arr[2581] : arr[2580];
wire r1_1292;
assign r1_1292 = in[0]? arr[2583] : arr[2582];
wire r1_1293;
assign r1_1293 = in[0]? arr[2585] : arr[2584];
wire r1_1294;
assign r1_1294 = in[0]? arr[2587] : arr[2586];
wire r1_1295;
assign r1_1295 = in[0]? arr[2589] : arr[2588];
wire r1_1296;
assign r1_1296 = in[0]? arr[2591] : arr[2590];
wire r1_1297;
assign r1_1297 = in[0]? arr[2593] : arr[2592];
wire r1_1298;
assign r1_1298 = in[0]? arr[2595] : arr[2594];
wire r1_1299;
assign r1_1299 = in[0]? arr[2597] : arr[2596];
wire r1_1300;
assign r1_1300 = in[0]? arr[2599] : arr[2598];
wire r1_1301;
assign r1_1301 = in[0]? arr[2601] : arr[2600];
wire r1_1302;
assign r1_1302 = in[0]? arr[2603] : arr[2602];
wire r1_1303;
assign r1_1303 = in[0]? arr[2605] : arr[2604];
wire r1_1304;
assign r1_1304 = in[0]? arr[2607] : arr[2606];
wire r1_1305;
assign r1_1305 = in[0]? arr[2609] : arr[2608];
wire r1_1306;
assign r1_1306 = in[0]? arr[2611] : arr[2610];
wire r1_1307;
assign r1_1307 = in[0]? arr[2613] : arr[2612];
wire r1_1308;
assign r1_1308 = in[0]? arr[2615] : arr[2614];
wire r1_1309;
assign r1_1309 = in[0]? arr[2617] : arr[2616];
wire r1_1310;
assign r1_1310 = in[0]? arr[2619] : arr[2618];
wire r1_1311;
assign r1_1311 = in[0]? arr[2621] : arr[2620];
wire r1_1312;
assign r1_1312 = in[0]? arr[2623] : arr[2622];
wire r1_1313;
assign r1_1313 = in[0]? arr[2625] : arr[2624];
wire r1_1314;
assign r1_1314 = in[0]? arr[2627] : arr[2626];
wire r1_1315;
assign r1_1315 = in[0]? arr[2629] : arr[2628];
wire r1_1316;
assign r1_1316 = in[0]? arr[2631] : arr[2630];
wire r1_1317;
assign r1_1317 = in[0]? arr[2633] : arr[2632];
wire r1_1318;
assign r1_1318 = in[0]? arr[2635] : arr[2634];
wire r1_1319;
assign r1_1319 = in[0]? arr[2637] : arr[2636];
wire r1_1320;
assign r1_1320 = in[0]? arr[2639] : arr[2638];
wire r1_1321;
assign r1_1321 = in[0]? arr[2641] : arr[2640];
wire r1_1322;
assign r1_1322 = in[0]? arr[2643] : arr[2642];
wire r1_1323;
assign r1_1323 = in[0]? arr[2645] : arr[2644];
wire r1_1324;
assign r1_1324 = in[0]? arr[2647] : arr[2646];
wire r1_1325;
assign r1_1325 = in[0]? arr[2649] : arr[2648];
wire r1_1326;
assign r1_1326 = in[0]? arr[2651] : arr[2650];
wire r1_1327;
assign r1_1327 = in[0]? arr[2653] : arr[2652];
wire r1_1328;
assign r1_1328 = in[0]? arr[2655] : arr[2654];
wire r1_1329;
assign r1_1329 = in[0]? arr[2657] : arr[2656];
wire r1_1330;
assign r1_1330 = in[0]? arr[2659] : arr[2658];
wire r1_1331;
assign r1_1331 = in[0]? arr[2661] : arr[2660];
wire r1_1332;
assign r1_1332 = in[0]? arr[2663] : arr[2662];
wire r1_1333;
assign r1_1333 = in[0]? arr[2665] : arr[2664];
wire r1_1334;
assign r1_1334 = in[0]? arr[2667] : arr[2666];
wire r1_1335;
assign r1_1335 = in[0]? arr[2669] : arr[2668];
wire r1_1336;
assign r1_1336 = in[0]? arr[2671] : arr[2670];
wire r1_1337;
assign r1_1337 = in[0]? arr[2673] : arr[2672];
wire r1_1338;
assign r1_1338 = in[0]? arr[2675] : arr[2674];
wire r1_1339;
assign r1_1339 = in[0]? arr[2677] : arr[2676];
wire r1_1340;
assign r1_1340 = in[0]? arr[2679] : arr[2678];
wire r1_1341;
assign r1_1341 = in[0]? arr[2681] : arr[2680];
wire r1_1342;
assign r1_1342 = in[0]? arr[2683] : arr[2682];
wire r1_1343;
assign r1_1343 = in[0]? arr[2685] : arr[2684];
wire r1_1344;
assign r1_1344 = in[0]? arr[2687] : arr[2686];
wire r1_1345;
assign r1_1345 = in[0]? arr[2689] : arr[2688];
wire r1_1346;
assign r1_1346 = in[0]? arr[2691] : arr[2690];
wire r1_1347;
assign r1_1347 = in[0]? arr[2693] : arr[2692];
wire r1_1348;
assign r1_1348 = in[0]? arr[2695] : arr[2694];
wire r1_1349;
assign r1_1349 = in[0]? arr[2697] : arr[2696];
wire r1_1350;
assign r1_1350 = in[0]? arr[2699] : arr[2698];
wire r1_1351;
assign r1_1351 = in[0]? arr[2701] : arr[2700];
wire r1_1352;
assign r1_1352 = in[0]? arr[2703] : arr[2702];
wire r1_1353;
assign r1_1353 = in[0]? arr[2705] : arr[2704];
wire r1_1354;
assign r1_1354 = in[0]? arr[2707] : arr[2706];
wire r1_1355;
assign r1_1355 = in[0]? arr[2709] : arr[2708];
wire r1_1356;
assign r1_1356 = in[0]? arr[2711] : arr[2710];
wire r1_1357;
assign r1_1357 = in[0]? arr[2713] : arr[2712];
wire r1_1358;
assign r1_1358 = in[0]? arr[2715] : arr[2714];
wire r1_1359;
assign r1_1359 = in[0]? arr[2717] : arr[2716];
wire r1_1360;
assign r1_1360 = in[0]? arr[2719] : arr[2718];
wire r1_1361;
assign r1_1361 = in[0]? arr[2721] : arr[2720];
wire r1_1362;
assign r1_1362 = in[0]? arr[2723] : arr[2722];
wire r1_1363;
assign r1_1363 = in[0]? arr[2725] : arr[2724];
wire r1_1364;
assign r1_1364 = in[0]? arr[2727] : arr[2726];
wire r1_1365;
assign r1_1365 = in[0]? arr[2729] : arr[2728];
wire r1_1366;
assign r1_1366 = in[0]? arr[2731] : arr[2730];
wire r1_1367;
assign r1_1367 = in[0]? arr[2733] : arr[2732];
wire r1_1368;
assign r1_1368 = in[0]? arr[2735] : arr[2734];
wire r1_1369;
assign r1_1369 = in[0]? arr[2737] : arr[2736];
wire r1_1370;
assign r1_1370 = in[0]? arr[2739] : arr[2738];
wire r1_1371;
assign r1_1371 = in[0]? arr[2741] : arr[2740];
wire r1_1372;
assign r1_1372 = in[0]? arr[2743] : arr[2742];
wire r1_1373;
assign r1_1373 = in[0]? arr[2745] : arr[2744];
wire r1_1374;
assign r1_1374 = in[0]? arr[2747] : arr[2746];
wire r1_1375;
assign r1_1375 = in[0]? arr[2749] : arr[2748];
wire r1_1376;
assign r1_1376 = in[0]? arr[2751] : arr[2750];
wire r1_1377;
assign r1_1377 = in[0]? arr[2753] : arr[2752];
wire r1_1378;
assign r1_1378 = in[0]? arr[2755] : arr[2754];
wire r1_1379;
assign r1_1379 = in[0]? arr[2757] : arr[2756];
wire r1_1380;
assign r1_1380 = in[0]? arr[2759] : arr[2758];
wire r1_1381;
assign r1_1381 = in[0]? arr[2761] : arr[2760];
wire r1_1382;
assign r1_1382 = in[0]? arr[2763] : arr[2762];
wire r1_1383;
assign r1_1383 = in[0]? arr[2765] : arr[2764];
wire r1_1384;
assign r1_1384 = in[0]? arr[2767] : arr[2766];
wire r1_1385;
assign r1_1385 = in[0]? arr[2769] : arr[2768];
wire r1_1386;
assign r1_1386 = in[0]? arr[2771] : arr[2770];
wire r1_1387;
assign r1_1387 = in[0]? arr[2773] : arr[2772];
wire r1_1388;
assign r1_1388 = in[0]? arr[2775] : arr[2774];
wire r1_1389;
assign r1_1389 = in[0]? arr[2777] : arr[2776];
wire r1_1390;
assign r1_1390 = in[0]? arr[2779] : arr[2778];
wire r1_1391;
assign r1_1391 = in[0]? arr[2781] : arr[2780];
wire r1_1392;
assign r1_1392 = in[0]? arr[2783] : arr[2782];
wire r1_1393;
assign r1_1393 = in[0]? arr[2785] : arr[2784];
wire r1_1394;
assign r1_1394 = in[0]? arr[2787] : arr[2786];
wire r1_1395;
assign r1_1395 = in[0]? arr[2789] : arr[2788];
wire r1_1396;
assign r1_1396 = in[0]? arr[2791] : arr[2790];
wire r1_1397;
assign r1_1397 = in[0]? arr[2793] : arr[2792];
wire r1_1398;
assign r1_1398 = in[0]? arr[2795] : arr[2794];
wire r1_1399;
assign r1_1399 = in[0]? arr[2797] : arr[2796];
wire r1_1400;
assign r1_1400 = in[0]? arr[2799] : arr[2798];
wire r1_1401;
assign r1_1401 = in[0]? arr[2801] : arr[2800];
wire r1_1402;
assign r1_1402 = in[0]? arr[2803] : arr[2802];
wire r1_1403;
assign r1_1403 = in[0]? arr[2805] : arr[2804];
wire r1_1404;
assign r1_1404 = in[0]? arr[2807] : arr[2806];
wire r1_1405;
assign r1_1405 = in[0]? arr[2809] : arr[2808];
wire r1_1406;
assign r1_1406 = in[0]? arr[2811] : arr[2810];
wire r1_1407;
assign r1_1407 = in[0]? arr[2813] : arr[2812];
wire r1_1408;
assign r1_1408 = in[0]? arr[2815] : arr[2814];
wire r1_1409;
assign r1_1409 = in[0]? arr[2817] : arr[2816];
wire r1_1410;
assign r1_1410 = in[0]? arr[2819] : arr[2818];
wire r1_1411;
assign r1_1411 = in[0]? arr[2821] : arr[2820];
wire r1_1412;
assign r1_1412 = in[0]? arr[2823] : arr[2822];
wire r1_1413;
assign r1_1413 = in[0]? arr[2825] : arr[2824];
wire r1_1414;
assign r1_1414 = in[0]? arr[2827] : arr[2826];
wire r1_1415;
assign r1_1415 = in[0]? arr[2829] : arr[2828];
wire r1_1416;
assign r1_1416 = in[0]? arr[2831] : arr[2830];
wire r1_1417;
assign r1_1417 = in[0]? arr[2833] : arr[2832];
wire r1_1418;
assign r1_1418 = in[0]? arr[2835] : arr[2834];
wire r1_1419;
assign r1_1419 = in[0]? arr[2837] : arr[2836];
wire r1_1420;
assign r1_1420 = in[0]? arr[2839] : arr[2838];
wire r1_1421;
assign r1_1421 = in[0]? arr[2841] : arr[2840];
wire r1_1422;
assign r1_1422 = in[0]? arr[2843] : arr[2842];
wire r1_1423;
assign r1_1423 = in[0]? arr[2845] : arr[2844];
wire r1_1424;
assign r1_1424 = in[0]? arr[2847] : arr[2846];
wire r1_1425;
assign r1_1425 = in[0]? arr[2849] : arr[2848];
wire r1_1426;
assign r1_1426 = in[0]? arr[2851] : arr[2850];
wire r1_1427;
assign r1_1427 = in[0]? arr[2853] : arr[2852];
wire r1_1428;
assign r1_1428 = in[0]? arr[2855] : arr[2854];
wire r1_1429;
assign r1_1429 = in[0]? arr[2857] : arr[2856];
wire r1_1430;
assign r1_1430 = in[0]? arr[2859] : arr[2858];
wire r1_1431;
assign r1_1431 = in[0]? arr[2861] : arr[2860];
wire r1_1432;
assign r1_1432 = in[0]? arr[2863] : arr[2862];
wire r1_1433;
assign r1_1433 = in[0]? arr[2865] : arr[2864];
wire r1_1434;
assign r1_1434 = in[0]? arr[2867] : arr[2866];
wire r1_1435;
assign r1_1435 = in[0]? arr[2869] : arr[2868];
wire r1_1436;
assign r1_1436 = in[0]? arr[2871] : arr[2870];
wire r1_1437;
assign r1_1437 = in[0]? arr[2873] : arr[2872];
wire r1_1438;
assign r1_1438 = in[0]? arr[2875] : arr[2874];
wire r1_1439;
assign r1_1439 = in[0]? arr[2877] : arr[2876];
wire r1_1440;
assign r1_1440 = in[0]? arr[2879] : arr[2878];
wire r1_1441;
assign r1_1441 = in[0]? arr[2881] : arr[2880];
wire r1_1442;
assign r1_1442 = in[0]? arr[2883] : arr[2882];
wire r1_1443;
assign r1_1443 = in[0]? arr[2885] : arr[2884];
wire r1_1444;
assign r1_1444 = in[0]? arr[2887] : arr[2886];
wire r1_1445;
assign r1_1445 = in[0]? arr[2889] : arr[2888];
wire r1_1446;
assign r1_1446 = in[0]? arr[2891] : arr[2890];
wire r1_1447;
assign r1_1447 = in[0]? arr[2893] : arr[2892];
wire r1_1448;
assign r1_1448 = in[0]? arr[2895] : arr[2894];
wire r1_1449;
assign r1_1449 = in[0]? arr[2897] : arr[2896];
wire r1_1450;
assign r1_1450 = in[0]? arr[2899] : arr[2898];
wire r1_1451;
assign r1_1451 = in[0]? arr[2901] : arr[2900];
wire r1_1452;
assign r1_1452 = in[0]? arr[2903] : arr[2902];
wire r1_1453;
assign r1_1453 = in[0]? arr[2905] : arr[2904];
wire r1_1454;
assign r1_1454 = in[0]? arr[2907] : arr[2906];
wire r1_1455;
assign r1_1455 = in[0]? arr[2909] : arr[2908];
wire r1_1456;
assign r1_1456 = in[0]? arr[2911] : arr[2910];
wire r1_1457;
assign r1_1457 = in[0]? arr[2913] : arr[2912];
wire r1_1458;
assign r1_1458 = in[0]? arr[2915] : arr[2914];
wire r1_1459;
assign r1_1459 = in[0]? arr[2917] : arr[2916];
wire r1_1460;
assign r1_1460 = in[0]? arr[2919] : arr[2918];
wire r1_1461;
assign r1_1461 = in[0]? arr[2921] : arr[2920];
wire r1_1462;
assign r1_1462 = in[0]? arr[2923] : arr[2922];
wire r1_1463;
assign r1_1463 = in[0]? arr[2925] : arr[2924];
wire r1_1464;
assign r1_1464 = in[0]? arr[2927] : arr[2926];
wire r1_1465;
assign r1_1465 = in[0]? arr[2929] : arr[2928];
wire r1_1466;
assign r1_1466 = in[0]? arr[2931] : arr[2930];
wire r1_1467;
assign r1_1467 = in[0]? arr[2933] : arr[2932];
wire r1_1468;
assign r1_1468 = in[0]? arr[2935] : arr[2934];
wire r1_1469;
assign r1_1469 = in[0]? arr[2937] : arr[2936];
wire r1_1470;
assign r1_1470 = in[0]? arr[2939] : arr[2938];
wire r1_1471;
assign r1_1471 = in[0]? arr[2941] : arr[2940];
wire r1_1472;
assign r1_1472 = in[0]? arr[2943] : arr[2942];
wire r1_1473;
assign r1_1473 = in[0]? arr[2945] : arr[2944];
wire r1_1474;
assign r1_1474 = in[0]? arr[2947] : arr[2946];
wire r1_1475;
assign r1_1475 = in[0]? arr[2949] : arr[2948];
wire r1_1476;
assign r1_1476 = in[0]? arr[2951] : arr[2950];
wire r1_1477;
assign r1_1477 = in[0]? arr[2953] : arr[2952];
wire r1_1478;
assign r1_1478 = in[0]? arr[2955] : arr[2954];
wire r1_1479;
assign r1_1479 = in[0]? arr[2957] : arr[2956];
wire r1_1480;
assign r1_1480 = in[0]? arr[2959] : arr[2958];
wire r1_1481;
assign r1_1481 = in[0]? arr[2961] : arr[2960];
wire r1_1482;
assign r1_1482 = in[0]? arr[2963] : arr[2962];
wire r1_1483;
assign r1_1483 = in[0]? arr[2965] : arr[2964];
wire r1_1484;
assign r1_1484 = in[0]? arr[2967] : arr[2966];
wire r1_1485;
assign r1_1485 = in[0]? arr[2969] : arr[2968];
wire r1_1486;
assign r1_1486 = in[0]? arr[2971] : arr[2970];
wire r1_1487;
assign r1_1487 = in[0]? arr[2973] : arr[2972];
wire r1_1488;
assign r1_1488 = in[0]? arr[2975] : arr[2974];
wire r1_1489;
assign r1_1489 = in[0]? arr[2977] : arr[2976];
wire r1_1490;
assign r1_1490 = in[0]? arr[2979] : arr[2978];
wire r1_1491;
assign r1_1491 = in[0]? arr[2981] : arr[2980];
wire r1_1492;
assign r1_1492 = in[0]? arr[2983] : arr[2982];
wire r1_1493;
assign r1_1493 = in[0]? arr[2985] : arr[2984];
wire r1_1494;
assign r1_1494 = in[0]? arr[2987] : arr[2986];
wire r1_1495;
assign r1_1495 = in[0]? arr[2989] : arr[2988];
wire r1_1496;
assign r1_1496 = in[0]? arr[2991] : arr[2990];
wire r1_1497;
assign r1_1497 = in[0]? arr[2993] : arr[2992];
wire r1_1498;
assign r1_1498 = in[0]? arr[2995] : arr[2994];
wire r1_1499;
assign r1_1499 = in[0]? arr[2997] : arr[2996];
wire r1_1500;
assign r1_1500 = in[0]? arr[2999] : arr[2998];
wire r1_1501;
assign r1_1501 = in[0]? arr[3001] : arr[3000];
wire r1_1502;
assign r1_1502 = in[0]? arr[3003] : arr[3002];
wire r1_1503;
assign r1_1503 = in[0]? arr[3005] : arr[3004];
wire r1_1504;
assign r1_1504 = in[0]? arr[3007] : arr[3006];
wire r1_1505;
assign r1_1505 = in[0]? arr[3009] : arr[3008];
wire r1_1506;
assign r1_1506 = in[0]? arr[3011] : arr[3010];
wire r1_1507;
assign r1_1507 = in[0]? arr[3013] : arr[3012];
wire r1_1508;
assign r1_1508 = in[0]? arr[3015] : arr[3014];
wire r1_1509;
assign r1_1509 = in[0]? arr[3017] : arr[3016];
wire r1_1510;
assign r1_1510 = in[0]? arr[3019] : arr[3018];
wire r1_1511;
assign r1_1511 = in[0]? arr[3021] : arr[3020];
wire r1_1512;
assign r1_1512 = in[0]? arr[3023] : arr[3022];
wire r1_1513;
assign r1_1513 = in[0]? arr[3025] : arr[3024];
wire r1_1514;
assign r1_1514 = in[0]? arr[3027] : arr[3026];
wire r1_1515;
assign r1_1515 = in[0]? arr[3029] : arr[3028];
wire r1_1516;
assign r1_1516 = in[0]? arr[3031] : arr[3030];
wire r1_1517;
assign r1_1517 = in[0]? arr[3033] : arr[3032];
wire r1_1518;
assign r1_1518 = in[0]? arr[3035] : arr[3034];
wire r1_1519;
assign r1_1519 = in[0]? arr[3037] : arr[3036];
wire r1_1520;
assign r1_1520 = in[0]? arr[3039] : arr[3038];
wire r1_1521;
assign r1_1521 = in[0]? arr[3041] : arr[3040];
wire r1_1522;
assign r1_1522 = in[0]? arr[3043] : arr[3042];
wire r1_1523;
assign r1_1523 = in[0]? arr[3045] : arr[3044];
wire r1_1524;
assign r1_1524 = in[0]? arr[3047] : arr[3046];
wire r1_1525;
assign r1_1525 = in[0]? arr[3049] : arr[3048];
wire r1_1526;
assign r1_1526 = in[0]? arr[3051] : arr[3050];
wire r1_1527;
assign r1_1527 = in[0]? arr[3053] : arr[3052];
wire r1_1528;
assign r1_1528 = in[0]? arr[3055] : arr[3054];
wire r1_1529;
assign r1_1529 = in[0]? arr[3057] : arr[3056];
wire r1_1530;
assign r1_1530 = in[0]? arr[3059] : arr[3058];
wire r1_1531;
assign r1_1531 = in[0]? arr[3061] : arr[3060];
wire r1_1532;
assign r1_1532 = in[0]? arr[3063] : arr[3062];
wire r1_1533;
assign r1_1533 = in[0]? arr[3065] : arr[3064];
wire r1_1534;
assign r1_1534 = in[0]? arr[3067] : arr[3066];
wire r1_1535;
assign r1_1535 = in[0]? arr[3069] : arr[3068];
wire r1_1536;
assign r1_1536 = in[0]? arr[3071] : arr[3070];
wire r1_1537;
assign r1_1537 = in[0]? arr[3073] : arr[3072];
wire r1_1538;
assign r1_1538 = in[0]? arr[3075] : arr[3074];
wire r1_1539;
assign r1_1539 = in[0]? arr[3077] : arr[3076];
wire r1_1540;
assign r1_1540 = in[0]? arr[3079] : arr[3078];
wire r1_1541;
assign r1_1541 = in[0]? arr[3081] : arr[3080];
wire r1_1542;
assign r1_1542 = in[0]? arr[3083] : arr[3082];
wire r1_1543;
assign r1_1543 = in[0]? arr[3085] : arr[3084];
wire r1_1544;
assign r1_1544 = in[0]? arr[3087] : arr[3086];
wire r1_1545;
assign r1_1545 = in[0]? arr[3089] : arr[3088];
wire r1_1546;
assign r1_1546 = in[0]? arr[3091] : arr[3090];
wire r1_1547;
assign r1_1547 = in[0]? arr[3093] : arr[3092];
wire r1_1548;
assign r1_1548 = in[0]? arr[3095] : arr[3094];
wire r1_1549;
assign r1_1549 = in[0]? arr[3097] : arr[3096];
wire r1_1550;
assign r1_1550 = in[0]? arr[3099] : arr[3098];
wire r1_1551;
assign r1_1551 = in[0]? arr[3101] : arr[3100];
wire r1_1552;
assign r1_1552 = in[0]? arr[3103] : arr[3102];
wire r1_1553;
assign r1_1553 = in[0]? arr[3105] : arr[3104];
wire r1_1554;
assign r1_1554 = in[0]? arr[3107] : arr[3106];
wire r1_1555;
assign r1_1555 = in[0]? arr[3109] : arr[3108];
wire r1_1556;
assign r1_1556 = in[0]? arr[3111] : arr[3110];
wire r1_1557;
assign r1_1557 = in[0]? arr[3113] : arr[3112];
wire r1_1558;
assign r1_1558 = in[0]? arr[3115] : arr[3114];
wire r1_1559;
assign r1_1559 = in[0]? arr[3117] : arr[3116];
wire r1_1560;
assign r1_1560 = in[0]? arr[3119] : arr[3118];
wire r1_1561;
assign r1_1561 = in[0]? arr[3121] : arr[3120];
wire r1_1562;
assign r1_1562 = in[0]? arr[3123] : arr[3122];
wire r1_1563;
assign r1_1563 = in[0]? arr[3125] : arr[3124];
wire r1_1564;
assign r1_1564 = in[0]? arr[3127] : arr[3126];
wire r1_1565;
assign r1_1565 = in[0]? arr[3129] : arr[3128];
wire r1_1566;
assign r1_1566 = in[0]? arr[3131] : arr[3130];
wire r1_1567;
assign r1_1567 = in[0]? arr[3133] : arr[3132];
wire r1_1568;
assign r1_1568 = in[0]? arr[3135] : arr[3134];
wire r1_1569;
assign r1_1569 = in[0]? arr[3137] : arr[3136];
wire r1_1570;
assign r1_1570 = in[0]? arr[3139] : arr[3138];
wire r1_1571;
assign r1_1571 = in[0]? arr[3141] : arr[3140];
wire r1_1572;
assign r1_1572 = in[0]? arr[3143] : arr[3142];
wire r1_1573;
assign r1_1573 = in[0]? arr[3145] : arr[3144];
wire r1_1574;
assign r1_1574 = in[0]? arr[3147] : arr[3146];
wire r1_1575;
assign r1_1575 = in[0]? arr[3149] : arr[3148];
wire r1_1576;
assign r1_1576 = in[0]? arr[3151] : arr[3150];
wire r1_1577;
assign r1_1577 = in[0]? arr[3153] : arr[3152];
wire r1_1578;
assign r1_1578 = in[0]? arr[3155] : arr[3154];
wire r1_1579;
assign r1_1579 = in[0]? arr[3157] : arr[3156];
wire r1_1580;
assign r1_1580 = in[0]? arr[3159] : arr[3158];
wire r1_1581;
assign r1_1581 = in[0]? arr[3161] : arr[3160];
wire r1_1582;
assign r1_1582 = in[0]? arr[3163] : arr[3162];
wire r1_1583;
assign r1_1583 = in[0]? arr[3165] : arr[3164];
wire r1_1584;
assign r1_1584 = in[0]? arr[3167] : arr[3166];
wire r1_1585;
assign r1_1585 = in[0]? arr[3169] : arr[3168];
wire r1_1586;
assign r1_1586 = in[0]? arr[3171] : arr[3170];
wire r1_1587;
assign r1_1587 = in[0]? arr[3173] : arr[3172];
wire r1_1588;
assign r1_1588 = in[0]? arr[3175] : arr[3174];
wire r1_1589;
assign r1_1589 = in[0]? arr[3177] : arr[3176];
wire r1_1590;
assign r1_1590 = in[0]? arr[3179] : arr[3178];
wire r1_1591;
assign r1_1591 = in[0]? arr[3181] : arr[3180];
wire r1_1592;
assign r1_1592 = in[0]? arr[3183] : arr[3182];
wire r1_1593;
assign r1_1593 = in[0]? arr[3185] : arr[3184];
wire r1_1594;
assign r1_1594 = in[0]? arr[3187] : arr[3186];
wire r1_1595;
assign r1_1595 = in[0]? arr[3189] : arr[3188];
wire r1_1596;
assign r1_1596 = in[0]? arr[3191] : arr[3190];
wire r1_1597;
assign r1_1597 = in[0]? arr[3193] : arr[3192];
wire r1_1598;
assign r1_1598 = in[0]? arr[3195] : arr[3194];
wire r1_1599;
assign r1_1599 = in[0]? arr[3197] : arr[3196];
wire r1_1600;
assign r1_1600 = in[0]? arr[3199] : arr[3198];
wire r1_1601;
assign r1_1601 = in[0]? arr[3201] : arr[3200];
wire r1_1602;
assign r1_1602 = in[0]? arr[3203] : arr[3202];
wire r1_1603;
assign r1_1603 = in[0]? arr[3205] : arr[3204];
wire r1_1604;
assign r1_1604 = in[0]? arr[3207] : arr[3206];
wire r1_1605;
assign r1_1605 = in[0]? arr[3209] : arr[3208];
wire r1_1606;
assign r1_1606 = in[0]? arr[3211] : arr[3210];
wire r1_1607;
assign r1_1607 = in[0]? arr[3213] : arr[3212];
wire r1_1608;
assign r1_1608 = in[0]? arr[3215] : arr[3214];
wire r1_1609;
assign r1_1609 = in[0]? arr[3217] : arr[3216];
wire r1_1610;
assign r1_1610 = in[0]? arr[3219] : arr[3218];
wire r1_1611;
assign r1_1611 = in[0]? arr[3221] : arr[3220];
wire r1_1612;
assign r1_1612 = in[0]? arr[3223] : arr[3222];
wire r1_1613;
assign r1_1613 = in[0]? arr[3225] : arr[3224];
wire r1_1614;
assign r1_1614 = in[0]? arr[3227] : arr[3226];
wire r1_1615;
assign r1_1615 = in[0]? arr[3229] : arr[3228];
wire r1_1616;
assign r1_1616 = in[0]? arr[3231] : arr[3230];
wire r1_1617;
assign r1_1617 = in[0]? arr[3233] : arr[3232];
wire r1_1618;
assign r1_1618 = in[0]? arr[3235] : arr[3234];
wire r1_1619;
assign r1_1619 = in[0]? arr[3237] : arr[3236];
wire r1_1620;
assign r1_1620 = in[0]? arr[3239] : arr[3238];
wire r1_1621;
assign r1_1621 = in[0]? arr[3241] : arr[3240];
wire r1_1622;
assign r1_1622 = in[0]? arr[3243] : arr[3242];
wire r1_1623;
assign r1_1623 = in[0]? arr[3245] : arr[3244];
wire r1_1624;
assign r1_1624 = in[0]? arr[3247] : arr[3246];
wire r1_1625;
assign r1_1625 = in[0]? arr[3249] : arr[3248];
wire r1_1626;
assign r1_1626 = in[0]? arr[3251] : arr[3250];
wire r1_1627;
assign r1_1627 = in[0]? arr[3253] : arr[3252];
wire r1_1628;
assign r1_1628 = in[0]? arr[3255] : arr[3254];
wire r1_1629;
assign r1_1629 = in[0]? arr[3257] : arr[3256];
wire r1_1630;
assign r1_1630 = in[0]? arr[3259] : arr[3258];
wire r1_1631;
assign r1_1631 = in[0]? arr[3261] : arr[3260];
wire r1_1632;
assign r1_1632 = in[0]? arr[3263] : arr[3262];
wire r1_1633;
assign r1_1633 = in[0]? arr[3265] : arr[3264];
wire r1_1634;
assign r1_1634 = in[0]? arr[3267] : arr[3266];
wire r1_1635;
assign r1_1635 = in[0]? arr[3269] : arr[3268];
wire r1_1636;
assign r1_1636 = in[0]? arr[3271] : arr[3270];
wire r1_1637;
assign r1_1637 = in[0]? arr[3273] : arr[3272];
wire r1_1638;
assign r1_1638 = in[0]? arr[3275] : arr[3274];
wire r1_1639;
assign r1_1639 = in[0]? arr[3277] : arr[3276];
wire r1_1640;
assign r1_1640 = in[0]? arr[3279] : arr[3278];
wire r1_1641;
assign r1_1641 = in[0]? arr[3281] : arr[3280];
wire r1_1642;
assign r1_1642 = in[0]? arr[3283] : arr[3282];
wire r1_1643;
assign r1_1643 = in[0]? arr[3285] : arr[3284];
wire r1_1644;
assign r1_1644 = in[0]? arr[3287] : arr[3286];
wire r1_1645;
assign r1_1645 = in[0]? arr[3289] : arr[3288];
wire r1_1646;
assign r1_1646 = in[0]? arr[3291] : arr[3290];
wire r1_1647;
assign r1_1647 = in[0]? arr[3293] : arr[3292];
wire r1_1648;
assign r1_1648 = in[0]? arr[3295] : arr[3294];
wire r1_1649;
assign r1_1649 = in[0]? arr[3297] : arr[3296];
wire r1_1650;
assign r1_1650 = in[0]? arr[3299] : arr[3298];
wire r1_1651;
assign r1_1651 = in[0]? arr[3301] : arr[3300];
wire r1_1652;
assign r1_1652 = in[0]? arr[3303] : arr[3302];
wire r1_1653;
assign r1_1653 = in[0]? arr[3305] : arr[3304];
wire r1_1654;
assign r1_1654 = in[0]? arr[3307] : arr[3306];
wire r1_1655;
assign r1_1655 = in[0]? arr[3309] : arr[3308];
wire r1_1656;
assign r1_1656 = in[0]? arr[3311] : arr[3310];
wire r1_1657;
assign r1_1657 = in[0]? arr[3313] : arr[3312];
wire r1_1658;
assign r1_1658 = in[0]? arr[3315] : arr[3314];
wire r1_1659;
assign r1_1659 = in[0]? arr[3317] : arr[3316];
wire r1_1660;
assign r1_1660 = in[0]? arr[3319] : arr[3318];
wire r1_1661;
assign r1_1661 = in[0]? arr[3321] : arr[3320];
wire r1_1662;
assign r1_1662 = in[0]? arr[3323] : arr[3322];
wire r1_1663;
assign r1_1663 = in[0]? arr[3325] : arr[3324];
wire r1_1664;
assign r1_1664 = in[0]? arr[3327] : arr[3326];
wire r1_1665;
assign r1_1665 = in[0]? arr[3329] : arr[3328];
wire r1_1666;
assign r1_1666 = in[0]? arr[3331] : arr[3330];
wire r1_1667;
assign r1_1667 = in[0]? arr[3333] : arr[3332];
wire r1_1668;
assign r1_1668 = in[0]? arr[3335] : arr[3334];
wire r1_1669;
assign r1_1669 = in[0]? arr[3337] : arr[3336];
wire r1_1670;
assign r1_1670 = in[0]? arr[3339] : arr[3338];
wire r1_1671;
assign r1_1671 = in[0]? arr[3341] : arr[3340];
wire r1_1672;
assign r1_1672 = in[0]? arr[3343] : arr[3342];
wire r1_1673;
assign r1_1673 = in[0]? arr[3345] : arr[3344];
wire r1_1674;
assign r1_1674 = in[0]? arr[3347] : arr[3346];
wire r1_1675;
assign r1_1675 = in[0]? arr[3349] : arr[3348];
wire r1_1676;
assign r1_1676 = in[0]? arr[3351] : arr[3350];
wire r1_1677;
assign r1_1677 = in[0]? arr[3353] : arr[3352];
wire r1_1678;
assign r1_1678 = in[0]? arr[3355] : arr[3354];
wire r1_1679;
assign r1_1679 = in[0]? arr[3357] : arr[3356];
wire r1_1680;
assign r1_1680 = in[0]? arr[3359] : arr[3358];
wire r1_1681;
assign r1_1681 = in[0]? arr[3361] : arr[3360];
wire r1_1682;
assign r1_1682 = in[0]? arr[3363] : arr[3362];
wire r1_1683;
assign r1_1683 = in[0]? arr[3365] : arr[3364];
wire r1_1684;
assign r1_1684 = in[0]? arr[3367] : arr[3366];
wire r1_1685;
assign r1_1685 = in[0]? arr[3369] : arr[3368];
wire r1_1686;
assign r1_1686 = in[0]? arr[3371] : arr[3370];
wire r1_1687;
assign r1_1687 = in[0]? arr[3373] : arr[3372];
wire r1_1688;
assign r1_1688 = in[0]? arr[3375] : arr[3374];
wire r1_1689;
assign r1_1689 = in[0]? arr[3377] : arr[3376];
wire r1_1690;
assign r1_1690 = in[0]? arr[3379] : arr[3378];
wire r1_1691;
assign r1_1691 = in[0]? arr[3381] : arr[3380];
wire r1_1692;
assign r1_1692 = in[0]? arr[3383] : arr[3382];
wire r1_1693;
assign r1_1693 = in[0]? arr[3385] : arr[3384];
wire r1_1694;
assign r1_1694 = in[0]? arr[3387] : arr[3386];
wire r1_1695;
assign r1_1695 = in[0]? arr[3389] : arr[3388];
wire r1_1696;
assign r1_1696 = in[0]? arr[3391] : arr[3390];
wire r1_1697;
assign r1_1697 = in[0]? arr[3393] : arr[3392];
wire r1_1698;
assign r1_1698 = in[0]? arr[3395] : arr[3394];
wire r1_1699;
assign r1_1699 = in[0]? arr[3397] : arr[3396];
wire r1_1700;
assign r1_1700 = in[0]? arr[3399] : arr[3398];
wire r1_1701;
assign r1_1701 = in[0]? arr[3401] : arr[3400];
wire r1_1702;
assign r1_1702 = in[0]? arr[3403] : arr[3402];
wire r1_1703;
assign r1_1703 = in[0]? arr[3405] : arr[3404];
wire r1_1704;
assign r1_1704 = in[0]? arr[3407] : arr[3406];
wire r1_1705;
assign r1_1705 = in[0]? arr[3409] : arr[3408];
wire r1_1706;
assign r1_1706 = in[0]? arr[3411] : arr[3410];
wire r1_1707;
assign r1_1707 = in[0]? arr[3413] : arr[3412];
wire r1_1708;
assign r1_1708 = in[0]? arr[3415] : arr[3414];
wire r1_1709;
assign r1_1709 = in[0]? arr[3417] : arr[3416];
wire r1_1710;
assign r1_1710 = in[0]? arr[3419] : arr[3418];
wire r1_1711;
assign r1_1711 = in[0]? arr[3421] : arr[3420];
wire r1_1712;
assign r1_1712 = in[0]? arr[3423] : arr[3422];
wire r1_1713;
assign r1_1713 = in[0]? arr[3425] : arr[3424];
wire r1_1714;
assign r1_1714 = in[0]? arr[3427] : arr[3426];
wire r1_1715;
assign r1_1715 = in[0]? arr[3429] : arr[3428];
wire r1_1716;
assign r1_1716 = in[0]? arr[3431] : arr[3430];
wire r1_1717;
assign r1_1717 = in[0]? arr[3433] : arr[3432];
wire r1_1718;
assign r1_1718 = in[0]? arr[3435] : arr[3434];
wire r1_1719;
assign r1_1719 = in[0]? arr[3437] : arr[3436];
wire r1_1720;
assign r1_1720 = in[0]? arr[3439] : arr[3438];
wire r1_1721;
assign r1_1721 = in[0]? arr[3441] : arr[3440];
wire r1_1722;
assign r1_1722 = in[0]? arr[3443] : arr[3442];
wire r1_1723;
assign r1_1723 = in[0]? arr[3445] : arr[3444];
wire r1_1724;
assign r1_1724 = in[0]? arr[3447] : arr[3446];
wire r1_1725;
assign r1_1725 = in[0]? arr[3449] : arr[3448];
wire r1_1726;
assign r1_1726 = in[0]? arr[3451] : arr[3450];
wire r1_1727;
assign r1_1727 = in[0]? arr[3453] : arr[3452];
wire r1_1728;
assign r1_1728 = in[0]? arr[3455] : arr[3454];
wire r1_1729;
assign r1_1729 = in[0]? arr[3457] : arr[3456];
wire r1_1730;
assign r1_1730 = in[0]? arr[3459] : arr[3458];
wire r1_1731;
assign r1_1731 = in[0]? arr[3461] : arr[3460];
wire r1_1732;
assign r1_1732 = in[0]? arr[3463] : arr[3462];
wire r1_1733;
assign r1_1733 = in[0]? arr[3465] : arr[3464];
wire r1_1734;
assign r1_1734 = in[0]? arr[3467] : arr[3466];
wire r1_1735;
assign r1_1735 = in[0]? arr[3469] : arr[3468];
wire r1_1736;
assign r1_1736 = in[0]? arr[3471] : arr[3470];
wire r1_1737;
assign r1_1737 = in[0]? arr[3473] : arr[3472];
wire r1_1738;
assign r1_1738 = in[0]? arr[3475] : arr[3474];
wire r1_1739;
assign r1_1739 = in[0]? arr[3477] : arr[3476];
wire r1_1740;
assign r1_1740 = in[0]? arr[3479] : arr[3478];
wire r1_1741;
assign r1_1741 = in[0]? arr[3481] : arr[3480];
wire r1_1742;
assign r1_1742 = in[0]? arr[3483] : arr[3482];
wire r1_1743;
assign r1_1743 = in[0]? arr[3485] : arr[3484];
wire r1_1744;
assign r1_1744 = in[0]? arr[3487] : arr[3486];
wire r1_1745;
assign r1_1745 = in[0]? arr[3489] : arr[3488];
wire r1_1746;
assign r1_1746 = in[0]? arr[3491] : arr[3490];
wire r1_1747;
assign r1_1747 = in[0]? arr[3493] : arr[3492];
wire r1_1748;
assign r1_1748 = in[0]? arr[3495] : arr[3494];
wire r1_1749;
assign r1_1749 = in[0]? arr[3497] : arr[3496];
wire r1_1750;
assign r1_1750 = in[0]? arr[3499] : arr[3498];
wire r1_1751;
assign r1_1751 = in[0]? arr[3501] : arr[3500];
wire r1_1752;
assign r1_1752 = in[0]? arr[3503] : arr[3502];
wire r1_1753;
assign r1_1753 = in[0]? arr[3505] : arr[3504];
wire r1_1754;
assign r1_1754 = in[0]? arr[3507] : arr[3506];
wire r1_1755;
assign r1_1755 = in[0]? arr[3509] : arr[3508];
wire r1_1756;
assign r1_1756 = in[0]? arr[3511] : arr[3510];
wire r1_1757;
assign r1_1757 = in[0]? arr[3513] : arr[3512];
wire r1_1758;
assign r1_1758 = in[0]? arr[3515] : arr[3514];
wire r1_1759;
assign r1_1759 = in[0]? arr[3517] : arr[3516];
wire r1_1760;
assign r1_1760 = in[0]? arr[3519] : arr[3518];
wire r1_1761;
assign r1_1761 = in[0]? arr[3521] : arr[3520];
wire r1_1762;
assign r1_1762 = in[0]? arr[3523] : arr[3522];
wire r1_1763;
assign r1_1763 = in[0]? arr[3525] : arr[3524];
wire r1_1764;
assign r1_1764 = in[0]? arr[3527] : arr[3526];
wire r1_1765;
assign r1_1765 = in[0]? arr[3529] : arr[3528];
wire r1_1766;
assign r1_1766 = in[0]? arr[3531] : arr[3530];
wire r1_1767;
assign r1_1767 = in[0]? arr[3533] : arr[3532];
wire r1_1768;
assign r1_1768 = in[0]? arr[3535] : arr[3534];
wire r1_1769;
assign r1_1769 = in[0]? arr[3537] : arr[3536];
wire r1_1770;
assign r1_1770 = in[0]? arr[3539] : arr[3538];
wire r1_1771;
assign r1_1771 = in[0]? arr[3541] : arr[3540];
wire r1_1772;
assign r1_1772 = in[0]? arr[3543] : arr[3542];
wire r1_1773;
assign r1_1773 = in[0]? arr[3545] : arr[3544];
wire r1_1774;
assign r1_1774 = in[0]? arr[3547] : arr[3546];
wire r1_1775;
assign r1_1775 = in[0]? arr[3549] : arr[3548];
wire r1_1776;
assign r1_1776 = in[0]? arr[3551] : arr[3550];
wire r1_1777;
assign r1_1777 = in[0]? arr[3553] : arr[3552];
wire r1_1778;
assign r1_1778 = in[0]? arr[3555] : arr[3554];
wire r1_1779;
assign r1_1779 = in[0]? arr[3557] : arr[3556];
wire r1_1780;
assign r1_1780 = in[0]? arr[3559] : arr[3558];
wire r1_1781;
assign r1_1781 = in[0]? arr[3561] : arr[3560];
wire r1_1782;
assign r1_1782 = in[0]? arr[3563] : arr[3562];
wire r1_1783;
assign r1_1783 = in[0]? arr[3565] : arr[3564];
wire r1_1784;
assign r1_1784 = in[0]? arr[3567] : arr[3566];
wire r1_1785;
assign r1_1785 = in[0]? arr[3569] : arr[3568];
wire r1_1786;
assign r1_1786 = in[0]? arr[3571] : arr[3570];
wire r1_1787;
assign r1_1787 = in[0]? arr[3573] : arr[3572];
wire r1_1788;
assign r1_1788 = in[0]? arr[3575] : arr[3574];
wire r1_1789;
assign r1_1789 = in[0]? arr[3577] : arr[3576];
wire r1_1790;
assign r1_1790 = in[0]? arr[3579] : arr[3578];
wire r1_1791;
assign r1_1791 = in[0]? arr[3581] : arr[3580];
wire r1_1792;
assign r1_1792 = in[0]? arr[3583] : arr[3582];
wire r1_1793;
assign r1_1793 = in[0]? arr[3585] : arr[3584];
wire r1_1794;
assign r1_1794 = in[0]? arr[3587] : arr[3586];
wire r1_1795;
assign r1_1795 = in[0]? arr[3589] : arr[3588];
wire r1_1796;
assign r1_1796 = in[0]? arr[3591] : arr[3590];
wire r1_1797;
assign r1_1797 = in[0]? arr[3593] : arr[3592];
wire r1_1798;
assign r1_1798 = in[0]? arr[3595] : arr[3594];
wire r1_1799;
assign r1_1799 = in[0]? arr[3597] : arr[3596];
wire r1_1800;
assign r1_1800 = in[0]? arr[3599] : arr[3598];
wire r1_1801;
assign r1_1801 = in[0]? arr[3601] : arr[3600];
wire r1_1802;
assign r1_1802 = in[0]? arr[3603] : arr[3602];
wire r1_1803;
assign r1_1803 = in[0]? arr[3605] : arr[3604];
wire r1_1804;
assign r1_1804 = in[0]? arr[3607] : arr[3606];
wire r1_1805;
assign r1_1805 = in[0]? arr[3609] : arr[3608];
wire r1_1806;
assign r1_1806 = in[0]? arr[3611] : arr[3610];
wire r1_1807;
assign r1_1807 = in[0]? arr[3613] : arr[3612];
wire r1_1808;
assign r1_1808 = in[0]? arr[3615] : arr[3614];
wire r1_1809;
assign r1_1809 = in[0]? arr[3617] : arr[3616];
wire r1_1810;
assign r1_1810 = in[0]? arr[3619] : arr[3618];
wire r1_1811;
assign r1_1811 = in[0]? arr[3621] : arr[3620];
wire r1_1812;
assign r1_1812 = in[0]? arr[3623] : arr[3622];
wire r1_1813;
assign r1_1813 = in[0]? arr[3625] : arr[3624];
wire r1_1814;
assign r1_1814 = in[0]? arr[3627] : arr[3626];
wire r1_1815;
assign r1_1815 = in[0]? arr[3629] : arr[3628];
wire r1_1816;
assign r1_1816 = in[0]? arr[3631] : arr[3630];
wire r1_1817;
assign r1_1817 = in[0]? arr[3633] : arr[3632];
wire r1_1818;
assign r1_1818 = in[0]? arr[3635] : arr[3634];
wire r1_1819;
assign r1_1819 = in[0]? arr[3637] : arr[3636];
wire r1_1820;
assign r1_1820 = in[0]? arr[3639] : arr[3638];
wire r1_1821;
assign r1_1821 = in[0]? arr[3641] : arr[3640];
wire r1_1822;
assign r1_1822 = in[0]? arr[3643] : arr[3642];
wire r1_1823;
assign r1_1823 = in[0]? arr[3645] : arr[3644];
wire r1_1824;
assign r1_1824 = in[0]? arr[3647] : arr[3646];
wire r1_1825;
assign r1_1825 = in[0]? arr[3649] : arr[3648];
wire r1_1826;
assign r1_1826 = in[0]? arr[3651] : arr[3650];
wire r1_1827;
assign r1_1827 = in[0]? arr[3653] : arr[3652];
wire r1_1828;
assign r1_1828 = in[0]? arr[3655] : arr[3654];
wire r1_1829;
assign r1_1829 = in[0]? arr[3657] : arr[3656];
wire r1_1830;
assign r1_1830 = in[0]? arr[3659] : arr[3658];
wire r1_1831;
assign r1_1831 = in[0]? arr[3661] : arr[3660];
wire r1_1832;
assign r1_1832 = in[0]? arr[3663] : arr[3662];
wire r1_1833;
assign r1_1833 = in[0]? arr[3665] : arr[3664];
wire r1_1834;
assign r1_1834 = in[0]? arr[3667] : arr[3666];
wire r1_1835;
assign r1_1835 = in[0]? arr[3669] : arr[3668];
wire r1_1836;
assign r1_1836 = in[0]? arr[3671] : arr[3670];
wire r1_1837;
assign r1_1837 = in[0]? arr[3673] : arr[3672];
wire r1_1838;
assign r1_1838 = in[0]? arr[3675] : arr[3674];
wire r1_1839;
assign r1_1839 = in[0]? arr[3677] : arr[3676];
wire r1_1840;
assign r1_1840 = in[0]? arr[3679] : arr[3678];
wire r1_1841;
assign r1_1841 = in[0]? arr[3681] : arr[3680];
wire r1_1842;
assign r1_1842 = in[0]? arr[3683] : arr[3682];
wire r1_1843;
assign r1_1843 = in[0]? arr[3685] : arr[3684];
wire r1_1844;
assign r1_1844 = in[0]? arr[3687] : arr[3686];
wire r1_1845;
assign r1_1845 = in[0]? arr[3689] : arr[3688];
wire r1_1846;
assign r1_1846 = in[0]? arr[3691] : arr[3690];
wire r1_1847;
assign r1_1847 = in[0]? arr[3693] : arr[3692];
wire r1_1848;
assign r1_1848 = in[0]? arr[3695] : arr[3694];
wire r1_1849;
assign r1_1849 = in[0]? arr[3697] : arr[3696];
wire r1_1850;
assign r1_1850 = in[0]? arr[3699] : arr[3698];
wire r1_1851;
assign r1_1851 = in[0]? arr[3701] : arr[3700];
wire r1_1852;
assign r1_1852 = in[0]? arr[3703] : arr[3702];
wire r1_1853;
assign r1_1853 = in[0]? arr[3705] : arr[3704];
wire r1_1854;
assign r1_1854 = in[0]? arr[3707] : arr[3706];
wire r1_1855;
assign r1_1855 = in[0]? arr[3709] : arr[3708];
wire r1_1856;
assign r1_1856 = in[0]? arr[3711] : arr[3710];
wire r1_1857;
assign r1_1857 = in[0]? arr[3713] : arr[3712];
wire r1_1858;
assign r1_1858 = in[0]? arr[3715] : arr[3714];
wire r1_1859;
assign r1_1859 = in[0]? arr[3717] : arr[3716];
wire r1_1860;
assign r1_1860 = in[0]? arr[3719] : arr[3718];
wire r1_1861;
assign r1_1861 = in[0]? arr[3721] : arr[3720];
wire r1_1862;
assign r1_1862 = in[0]? arr[3723] : arr[3722];
wire r1_1863;
assign r1_1863 = in[0]? arr[3725] : arr[3724];
wire r1_1864;
assign r1_1864 = in[0]? arr[3727] : arr[3726];
wire r1_1865;
assign r1_1865 = in[0]? arr[3729] : arr[3728];
wire r1_1866;
assign r1_1866 = in[0]? arr[3731] : arr[3730];
wire r1_1867;
assign r1_1867 = in[0]? arr[3733] : arr[3732];
wire r1_1868;
assign r1_1868 = in[0]? arr[3735] : arr[3734];
wire r1_1869;
assign r1_1869 = in[0]? arr[3737] : arr[3736];
wire r1_1870;
assign r1_1870 = in[0]? arr[3739] : arr[3738];
wire r1_1871;
assign r1_1871 = in[0]? arr[3741] : arr[3740];
wire r1_1872;
assign r1_1872 = in[0]? arr[3743] : arr[3742];
wire r1_1873;
assign r1_1873 = in[0]? arr[3745] : arr[3744];
wire r1_1874;
assign r1_1874 = in[0]? arr[3747] : arr[3746];
wire r1_1875;
assign r1_1875 = in[0]? arr[3749] : arr[3748];
wire r1_1876;
assign r1_1876 = in[0]? arr[3751] : arr[3750];
wire r1_1877;
assign r1_1877 = in[0]? arr[3753] : arr[3752];
wire r1_1878;
assign r1_1878 = in[0]? arr[3755] : arr[3754];
wire r1_1879;
assign r1_1879 = in[0]? arr[3757] : arr[3756];
wire r1_1880;
assign r1_1880 = in[0]? arr[3759] : arr[3758];
wire r1_1881;
assign r1_1881 = in[0]? arr[3761] : arr[3760];
wire r1_1882;
assign r1_1882 = in[0]? arr[3763] : arr[3762];
wire r1_1883;
assign r1_1883 = in[0]? arr[3765] : arr[3764];
wire r1_1884;
assign r1_1884 = in[0]? arr[3767] : arr[3766];
wire r1_1885;
assign r1_1885 = in[0]? arr[3769] : arr[3768];
wire r1_1886;
assign r1_1886 = in[0]? arr[3771] : arr[3770];
wire r1_1887;
assign r1_1887 = in[0]? arr[3773] : arr[3772];
wire r1_1888;
assign r1_1888 = in[0]? arr[3775] : arr[3774];
wire r1_1889;
assign r1_1889 = in[0]? arr[3777] : arr[3776];
wire r1_1890;
assign r1_1890 = in[0]? arr[3779] : arr[3778];
wire r1_1891;
assign r1_1891 = in[0]? arr[3781] : arr[3780];
wire r1_1892;
assign r1_1892 = in[0]? arr[3783] : arr[3782];
wire r1_1893;
assign r1_1893 = in[0]? arr[3785] : arr[3784];
wire r1_1894;
assign r1_1894 = in[0]? arr[3787] : arr[3786];
wire r1_1895;
assign r1_1895 = in[0]? arr[3789] : arr[3788];
wire r1_1896;
assign r1_1896 = in[0]? arr[3791] : arr[3790];
wire r1_1897;
assign r1_1897 = in[0]? arr[3793] : arr[3792];
wire r1_1898;
assign r1_1898 = in[0]? arr[3795] : arr[3794];
wire r1_1899;
assign r1_1899 = in[0]? arr[3797] : arr[3796];
wire r1_1900;
assign r1_1900 = in[0]? arr[3799] : arr[3798];
wire r1_1901;
assign r1_1901 = in[0]? arr[3801] : arr[3800];
wire r1_1902;
assign r1_1902 = in[0]? arr[3803] : arr[3802];
wire r1_1903;
assign r1_1903 = in[0]? arr[3805] : arr[3804];
wire r1_1904;
assign r1_1904 = in[0]? arr[3807] : arr[3806];
wire r1_1905;
assign r1_1905 = in[0]? arr[3809] : arr[3808];
wire r1_1906;
assign r1_1906 = in[0]? arr[3811] : arr[3810];
wire r1_1907;
assign r1_1907 = in[0]? arr[3813] : arr[3812];
wire r1_1908;
assign r1_1908 = in[0]? arr[3815] : arr[3814];
wire r1_1909;
assign r1_1909 = in[0]? arr[3817] : arr[3816];
wire r1_1910;
assign r1_1910 = in[0]? arr[3819] : arr[3818];
wire r1_1911;
assign r1_1911 = in[0]? arr[3821] : arr[3820];
wire r1_1912;
assign r1_1912 = in[0]? arr[3823] : arr[3822];
wire r1_1913;
assign r1_1913 = in[0]? arr[3825] : arr[3824];
wire r1_1914;
assign r1_1914 = in[0]? arr[3827] : arr[3826];
wire r1_1915;
assign r1_1915 = in[0]? arr[3829] : arr[3828];
wire r1_1916;
assign r1_1916 = in[0]? arr[3831] : arr[3830];
wire r1_1917;
assign r1_1917 = in[0]? arr[3833] : arr[3832];
wire r1_1918;
assign r1_1918 = in[0]? arr[3835] : arr[3834];
wire r1_1919;
assign r1_1919 = in[0]? arr[3837] : arr[3836];
wire r1_1920;
assign r1_1920 = in[0]? arr[3839] : arr[3838];
wire r1_1921;
assign r1_1921 = in[0]? arr[3841] : arr[3840];
wire r1_1922;
assign r1_1922 = in[0]? arr[3843] : arr[3842];
wire r1_1923;
assign r1_1923 = in[0]? arr[3845] : arr[3844];
wire r1_1924;
assign r1_1924 = in[0]? arr[3847] : arr[3846];
wire r1_1925;
assign r1_1925 = in[0]? arr[3849] : arr[3848];
wire r1_1926;
assign r1_1926 = in[0]? arr[3851] : arr[3850];
wire r1_1927;
assign r1_1927 = in[0]? arr[3853] : arr[3852];
wire r1_1928;
assign r1_1928 = in[0]? arr[3855] : arr[3854];
wire r1_1929;
assign r1_1929 = in[0]? arr[3857] : arr[3856];
wire r1_1930;
assign r1_1930 = in[0]? arr[3859] : arr[3858];
wire r1_1931;
assign r1_1931 = in[0]? arr[3861] : arr[3860];
wire r1_1932;
assign r1_1932 = in[0]? arr[3863] : arr[3862];
wire r1_1933;
assign r1_1933 = in[0]? arr[3865] : arr[3864];
wire r1_1934;
assign r1_1934 = in[0]? arr[3867] : arr[3866];
wire r1_1935;
assign r1_1935 = in[0]? arr[3869] : arr[3868];
wire r1_1936;
assign r1_1936 = in[0]? arr[3871] : arr[3870];
wire r1_1937;
assign r1_1937 = in[0]? arr[3873] : arr[3872];
wire r1_1938;
assign r1_1938 = in[0]? arr[3875] : arr[3874];
wire r1_1939;
assign r1_1939 = in[0]? arr[3877] : arr[3876];
wire r1_1940;
assign r1_1940 = in[0]? arr[3879] : arr[3878];
wire r1_1941;
assign r1_1941 = in[0]? arr[3881] : arr[3880];
wire r1_1942;
assign r1_1942 = in[0]? arr[3883] : arr[3882];
wire r1_1943;
assign r1_1943 = in[0]? arr[3885] : arr[3884];
wire r1_1944;
assign r1_1944 = in[0]? arr[3887] : arr[3886];
wire r1_1945;
assign r1_1945 = in[0]? arr[3889] : arr[3888];
wire r1_1946;
assign r1_1946 = in[0]? arr[3891] : arr[3890];
wire r1_1947;
assign r1_1947 = in[0]? arr[3893] : arr[3892];
wire r1_1948;
assign r1_1948 = in[0]? arr[3895] : arr[3894];
wire r1_1949;
assign r1_1949 = in[0]? arr[3897] : arr[3896];
wire r1_1950;
assign r1_1950 = in[0]? arr[3899] : arr[3898];
wire r1_1951;
assign r1_1951 = in[0]? arr[3901] : arr[3900];
wire r1_1952;
assign r1_1952 = in[0]? arr[3903] : arr[3902];
wire r1_1953;
assign r1_1953 = in[0]? arr[3905] : arr[3904];
wire r1_1954;
assign r1_1954 = in[0]? arr[3907] : arr[3906];
wire r1_1955;
assign r1_1955 = in[0]? arr[3909] : arr[3908];
wire r1_1956;
assign r1_1956 = in[0]? arr[3911] : arr[3910];
wire r1_1957;
assign r1_1957 = in[0]? arr[3913] : arr[3912];
wire r1_1958;
assign r1_1958 = in[0]? arr[3915] : arr[3914];
wire r1_1959;
assign r1_1959 = in[0]? arr[3917] : arr[3916];
wire r1_1960;
assign r1_1960 = in[0]? arr[3919] : arr[3918];
wire r1_1961;
assign r1_1961 = in[0]? arr[3921] : arr[3920];
wire r1_1962;
assign r1_1962 = in[0]? arr[3923] : arr[3922];
wire r1_1963;
assign r1_1963 = in[0]? arr[3925] : arr[3924];
wire r1_1964;
assign r1_1964 = in[0]? arr[3927] : arr[3926];
wire r1_1965;
assign r1_1965 = in[0]? arr[3929] : arr[3928];
wire r1_1966;
assign r1_1966 = in[0]? arr[3931] : arr[3930];
wire r1_1967;
assign r1_1967 = in[0]? arr[3933] : arr[3932];
wire r1_1968;
assign r1_1968 = in[0]? arr[3935] : arr[3934];
wire r1_1969;
assign r1_1969 = in[0]? arr[3937] : arr[3936];
wire r1_1970;
assign r1_1970 = in[0]? arr[3939] : arr[3938];
wire r1_1971;
assign r1_1971 = in[0]? arr[3941] : arr[3940];
wire r1_1972;
assign r1_1972 = in[0]? arr[3943] : arr[3942];
wire r1_1973;
assign r1_1973 = in[0]? arr[3945] : arr[3944];
wire r1_1974;
assign r1_1974 = in[0]? arr[3947] : arr[3946];
wire r1_1975;
assign r1_1975 = in[0]? arr[3949] : arr[3948];
wire r1_1976;
assign r1_1976 = in[0]? arr[3951] : arr[3950];
wire r1_1977;
assign r1_1977 = in[0]? arr[3953] : arr[3952];
wire r1_1978;
assign r1_1978 = in[0]? arr[3955] : arr[3954];
wire r1_1979;
assign r1_1979 = in[0]? arr[3957] : arr[3956];
wire r1_1980;
assign r1_1980 = in[0]? arr[3959] : arr[3958];
wire r1_1981;
assign r1_1981 = in[0]? arr[3961] : arr[3960];
wire r1_1982;
assign r1_1982 = in[0]? arr[3963] : arr[3962];
wire r1_1983;
assign r1_1983 = in[0]? arr[3965] : arr[3964];
wire r1_1984;
assign r1_1984 = in[0]? arr[3967] : arr[3966];
wire r1_1985;
assign r1_1985 = in[0]? arr[3969] : arr[3968];
wire r1_1986;
assign r1_1986 = in[0]? arr[3971] : arr[3970];
wire r1_1987;
assign r1_1987 = in[0]? arr[3973] : arr[3972];
wire r1_1988;
assign r1_1988 = in[0]? arr[3975] : arr[3974];
wire r1_1989;
assign r1_1989 = in[0]? arr[3977] : arr[3976];
wire r1_1990;
assign r1_1990 = in[0]? arr[3979] : arr[3978];
wire r1_1991;
assign r1_1991 = in[0]? arr[3981] : arr[3980];
wire r1_1992;
assign r1_1992 = in[0]? arr[3983] : arr[3982];
wire r1_1993;
assign r1_1993 = in[0]? arr[3985] : arr[3984];
wire r1_1994;
assign r1_1994 = in[0]? arr[3987] : arr[3986];
wire r1_1995;
assign r1_1995 = in[0]? arr[3989] : arr[3988];
wire r1_1996;
assign r1_1996 = in[0]? arr[3991] : arr[3990];
wire r1_1997;
assign r1_1997 = in[0]? arr[3993] : arr[3992];
wire r1_1998;
assign r1_1998 = in[0]? arr[3995] : arr[3994];
wire r1_1999;
assign r1_1999 = in[0]? arr[3997] : arr[3996];
wire r1_2000;
assign r1_2000 = in[0]? arr[3999] : arr[3998];
wire r1_2001;
assign r1_2001 = in[0]? arr[4001] : arr[4000];
wire r1_2002;
assign r1_2002 = in[0]? arr[4003] : arr[4002];
wire r1_2003;
assign r1_2003 = in[0]? arr[4005] : arr[4004];
wire r1_2004;
assign r1_2004 = in[0]? arr[4007] : arr[4006];
wire r1_2005;
assign r1_2005 = in[0]? arr[4009] : arr[4008];
wire r1_2006;
assign r1_2006 = in[0]? arr[4011] : arr[4010];
wire r1_2007;
assign r1_2007 = in[0]? arr[4013] : arr[4012];
wire r1_2008;
assign r1_2008 = in[0]? arr[4015] : arr[4014];
wire r1_2009;
assign r1_2009 = in[0]? arr[4017] : arr[4016];
wire r1_2010;
assign r1_2010 = in[0]? arr[4019] : arr[4018];
wire r1_2011;
assign r1_2011 = in[0]? arr[4021] : arr[4020];
wire r1_2012;
assign r1_2012 = in[0]? arr[4023] : arr[4022];
wire r1_2013;
assign r1_2013 = in[0]? arr[4025] : arr[4024];
wire r1_2014;
assign r1_2014 = in[0]? arr[4027] : arr[4026];
wire r1_2015;
assign r1_2015 = in[0]? arr[4029] : arr[4028];
wire r1_2016;
assign r1_2016 = in[0]? arr[4031] : arr[4030];
wire r1_2017;
assign r1_2017 = in[0]? arr[4033] : arr[4032];
wire r1_2018;
assign r1_2018 = in[0]? arr[4035] : arr[4034];
wire r1_2019;
assign r1_2019 = in[0]? arr[4037] : arr[4036];
wire r1_2020;
assign r1_2020 = in[0]? arr[4039] : arr[4038];
wire r1_2021;
assign r1_2021 = in[0]? arr[4041] : arr[4040];
wire r1_2022;
assign r1_2022 = in[0]? arr[4043] : arr[4042];
wire r1_2023;
assign r1_2023 = in[0]? arr[4045] : arr[4044];
wire r1_2024;
assign r1_2024 = in[0]? arr[4047] : arr[4046];
wire r1_2025;
assign r1_2025 = in[0]? arr[4049] : arr[4048];
wire r1_2026;
assign r1_2026 = in[0]? arr[4051] : arr[4050];
wire r1_2027;
assign r1_2027 = in[0]? arr[4053] : arr[4052];
wire r1_2028;
assign r1_2028 = in[0]? arr[4055] : arr[4054];
wire r1_2029;
assign r1_2029 = in[0]? arr[4057] : arr[4056];
wire r1_2030;
assign r1_2030 = in[0]? arr[4059] : arr[4058];
wire r1_2031;
assign r1_2031 = in[0]? arr[4061] : arr[4060];
wire r1_2032;
assign r1_2032 = in[0]? arr[4063] : arr[4062];
wire r1_2033;
assign r1_2033 = in[0]? arr[4065] : arr[4064];
wire r1_2034;
assign r1_2034 = in[0]? arr[4067] : arr[4066];
wire r1_2035;
assign r1_2035 = in[0]? arr[4069] : arr[4068];
wire r1_2036;
assign r1_2036 = in[0]? arr[4071] : arr[4070];
wire r1_2037;
assign r1_2037 = in[0]? arr[4073] : arr[4072];
wire r1_2038;
assign r1_2038 = in[0]? arr[4075] : arr[4074];
wire r1_2039;
assign r1_2039 = in[0]? arr[4077] : arr[4076];
wire r1_2040;
assign r1_2040 = in[0]? arr[4079] : arr[4078];
wire r1_2041;
assign r1_2041 = in[0]? arr[4081] : arr[4080];
wire r1_2042;
assign r1_2042 = in[0]? arr[4083] : arr[4082];
wire r1_2043;
assign r1_2043 = in[0]? arr[4085] : arr[4084];
wire r1_2044;
assign r1_2044 = in[0]? arr[4087] : arr[4086];
wire r1_2045;
assign r1_2045 = in[0]? arr[4089] : arr[4088];
wire r1_2046;
assign r1_2046 = in[0]? arr[4091] : arr[4090];
wire r1_2047;
assign r1_2047 = in[0]? arr[4093] : arr[4092];
wire r1_2048;
assign r1_2048 = in[0]? arr[4095] : arr[4094];
wire r1_2049;
assign r1_2049 = in[0]? arr[4097] : arr[4096];
wire r1_2050;
assign r1_2050 = in[0]? arr[4099] : arr[4098];
wire r1_2051;
assign r1_2051 = in[0]? arr[4101] : arr[4100];
wire r1_2052;
assign r1_2052 = in[0]? arr[4103] : arr[4102];
wire r1_2053;
assign r1_2053 = in[0]? arr[4105] : arr[4104];
wire r1_2054;
assign r1_2054 = in[0]? arr[4107] : arr[4106];
wire r1_2055;
assign r1_2055 = in[0]? arr[4109] : arr[4108];
wire r1_2056;
assign r1_2056 = in[0]? arr[4111] : arr[4110];
wire r1_2057;
assign r1_2057 = in[0]? arr[4113] : arr[4112];
wire r1_2058;
assign r1_2058 = in[0]? arr[4115] : arr[4114];
wire r1_2059;
assign r1_2059 = in[0]? arr[4117] : arr[4116];
wire r1_2060;
assign r1_2060 = in[0]? arr[4119] : arr[4118];
wire r1_2061;
assign r1_2061 = in[0]? arr[4121] : arr[4120];
wire r1_2062;
assign r1_2062 = in[0]? arr[4123] : arr[4122];
wire r1_2063;
assign r1_2063 = in[0]? arr[4125] : arr[4124];
wire r1_2064;
assign r1_2064 = in[0]? arr[4127] : arr[4126];
wire r1_2065;
assign r1_2065 = in[0]? arr[4129] : arr[4128];
wire r1_2066;
assign r1_2066 = in[0]? arr[4131] : arr[4130];
wire r1_2067;
assign r1_2067 = in[0]? arr[4133] : arr[4132];
wire r1_2068;
assign r1_2068 = in[0]? arr[4135] : arr[4134];
wire r1_2069;
assign r1_2069 = in[0]? arr[4137] : arr[4136];
wire r1_2070;
assign r1_2070 = in[0]? arr[4139] : arr[4138];
wire r1_2071;
assign r1_2071 = in[0]? arr[4141] : arr[4140];
wire r1_2072;
assign r1_2072 = in[0]? arr[4143] : arr[4142];
wire r1_2073;
assign r1_2073 = in[0]? arr[4145] : arr[4144];
wire r1_2074;
assign r1_2074 = in[0]? arr[4147] : arr[4146];
wire r1_2075;
assign r1_2075 = in[0]? arr[4149] : arr[4148];
wire r1_2076;
assign r1_2076 = in[0]? arr[4151] : arr[4150];
wire r1_2077;
assign r1_2077 = in[0]? arr[4153] : arr[4152];
wire r1_2078;
assign r1_2078 = in[0]? arr[4155] : arr[4154];
wire r1_2079;
assign r1_2079 = in[0]? arr[4157] : arr[4156];
wire r1_2080;
assign r1_2080 = in[0]? arr[4159] : arr[4158];
wire r1_2081;
assign r1_2081 = in[0]? arr[4161] : arr[4160];
wire r1_2082;
assign r1_2082 = in[0]? arr[4163] : arr[4162];
wire r1_2083;
assign r1_2083 = in[0]? arr[4165] : arr[4164];
wire r1_2084;
assign r1_2084 = in[0]? arr[4167] : arr[4166];
wire r1_2085;
assign r1_2085 = in[0]? arr[4169] : arr[4168];
wire r1_2086;
assign r1_2086 = in[0]? arr[4171] : arr[4170];
wire r1_2087;
assign r1_2087 = in[0]? arr[4173] : arr[4172];
wire r1_2088;
assign r1_2088 = in[0]? arr[4175] : arr[4174];
wire r1_2089;
assign r1_2089 = in[0]? arr[4177] : arr[4176];
wire r1_2090;
assign r1_2090 = in[0]? arr[4179] : arr[4178];
wire r1_2091;
assign r1_2091 = in[0]? arr[4181] : arr[4180];
wire r1_2092;
assign r1_2092 = in[0]? arr[4183] : arr[4182];
wire r1_2093;
assign r1_2093 = in[0]? arr[4185] : arr[4184];
wire r1_2094;
assign r1_2094 = in[0]? arr[4187] : arr[4186];
wire r1_2095;
assign r1_2095 = in[0]? arr[4189] : arr[4188];
wire r1_2096;
assign r1_2096 = in[0]? arr[4191] : arr[4190];
wire r1_2097;
assign r1_2097 = in[0]? arr[4193] : arr[4192];
wire r1_2098;
assign r1_2098 = in[0]? arr[4195] : arr[4194];
wire r1_2099;
assign r1_2099 = in[0]? arr[4197] : arr[4196];
wire r1_2100;
assign r1_2100 = in[0]? arr[4199] : arr[4198];
wire r1_2101;
assign r1_2101 = in[0]? arr[4201] : arr[4200];
wire r1_2102;
assign r1_2102 = in[0]? arr[4203] : arr[4202];
wire r1_2103;
assign r1_2103 = in[0]? arr[4205] : arr[4204];
wire r1_2104;
assign r1_2104 = in[0]? arr[4207] : arr[4206];
wire r1_2105;
assign r1_2105 = in[0]? arr[4209] : arr[4208];
wire r1_2106;
assign r1_2106 = in[0]? arr[4211] : arr[4210];
wire r1_2107;
assign r1_2107 = in[0]? arr[4213] : arr[4212];
wire r1_2108;
assign r1_2108 = in[0]? arr[4215] : arr[4214];
wire r1_2109;
assign r1_2109 = in[0]? arr[4217] : arr[4216];
wire r1_2110;
assign r1_2110 = in[0]? arr[4219] : arr[4218];
wire r1_2111;
assign r1_2111 = in[0]? arr[4221] : arr[4220];
wire r1_2112;
assign r1_2112 = in[0]? arr[4223] : arr[4222];
wire r1_2113;
assign r1_2113 = in[0]? arr[4225] : arr[4224];
wire r1_2114;
assign r1_2114 = in[0]? arr[4227] : arr[4226];
wire r1_2115;
assign r1_2115 = in[0]? arr[4229] : arr[4228];
wire r1_2116;
assign r1_2116 = in[0]? arr[4231] : arr[4230];
wire r1_2117;
assign r1_2117 = in[0]? arr[4233] : arr[4232];
wire r1_2118;
assign r1_2118 = in[0]? arr[4235] : arr[4234];
wire r1_2119;
assign r1_2119 = in[0]? arr[4237] : arr[4236];
wire r1_2120;
assign r1_2120 = in[0]? arr[4239] : arr[4238];
wire r1_2121;
assign r1_2121 = in[0]? arr[4241] : arr[4240];
wire r1_2122;
assign r1_2122 = in[0]? arr[4243] : arr[4242];
wire r1_2123;
assign r1_2123 = in[0]? arr[4245] : arr[4244];
wire r1_2124;
assign r1_2124 = in[0]? arr[4247] : arr[4246];
wire r1_2125;
assign r1_2125 = in[0]? arr[4249] : arr[4248];
wire r1_2126;
assign r1_2126 = in[0]? arr[4251] : arr[4250];
wire r1_2127;
assign r1_2127 = in[0]? arr[4253] : arr[4252];
wire r1_2128;
assign r1_2128 = in[0]? arr[4255] : arr[4254];
wire r1_2129;
assign r1_2129 = in[0]? arr[4257] : arr[4256];
wire r1_2130;
assign r1_2130 = in[0]? arr[4259] : arr[4258];
wire r1_2131;
assign r1_2131 = in[0]? arr[4261] : arr[4260];
wire r1_2132;
assign r1_2132 = in[0]? arr[4263] : arr[4262];
wire r1_2133;
assign r1_2133 = in[0]? arr[4265] : arr[4264];
wire r1_2134;
assign r1_2134 = in[0]? arr[4267] : arr[4266];
wire r1_2135;
assign r1_2135 = in[0]? arr[4269] : arr[4268];
wire r1_2136;
assign r1_2136 = in[0]? arr[4271] : arr[4270];
wire r1_2137;
assign r1_2137 = in[0]? arr[4273] : arr[4272];
wire r1_2138;
assign r1_2138 = in[0]? arr[4275] : arr[4274];
wire r1_2139;
assign r1_2139 = in[0]? arr[4277] : arr[4276];
wire r1_2140;
assign r1_2140 = in[0]? arr[4279] : arr[4278];
wire r1_2141;
assign r1_2141 = in[0]? arr[4281] : arr[4280];
wire r1_2142;
assign r1_2142 = in[0]? arr[4283] : arr[4282];
wire r1_2143;
assign r1_2143 = in[0]? arr[4285] : arr[4284];
wire r1_2144;
assign r1_2144 = in[0]? arr[4287] : arr[4286];
wire r1_2145;
assign r1_2145 = in[0]? arr[4289] : arr[4288];
wire r1_2146;
assign r1_2146 = in[0]? arr[4291] : arr[4290];
wire r1_2147;
assign r1_2147 = in[0]? arr[4293] : arr[4292];
wire r1_2148;
assign r1_2148 = in[0]? arr[4295] : arr[4294];
wire r1_2149;
assign r1_2149 = in[0]? arr[4297] : arr[4296];
wire r1_2150;
assign r1_2150 = in[0]? arr[4299] : arr[4298];
wire r1_2151;
assign r1_2151 = in[0]? arr[4301] : arr[4300];
wire r1_2152;
assign r1_2152 = in[0]? arr[4303] : arr[4302];
wire r1_2153;
assign r1_2153 = in[0]? arr[4305] : arr[4304];
wire r1_2154;
assign r1_2154 = in[0]? arr[4307] : arr[4306];
wire r1_2155;
assign r1_2155 = in[0]? arr[4309] : arr[4308];
wire r1_2156;
assign r1_2156 = in[0]? arr[4311] : arr[4310];
wire r1_2157;
assign r1_2157 = in[0]? arr[4313] : arr[4312];
wire r1_2158;
assign r1_2158 = in[0]? arr[4315] : arr[4314];
wire r1_2159;
assign r1_2159 = in[0]? arr[4317] : arr[4316];
wire r1_2160;
assign r1_2160 = in[0]? arr[4319] : arr[4318];
wire r1_2161;
assign r1_2161 = in[0]? arr[4321] : arr[4320];
wire r1_2162;
assign r1_2162 = in[0]? arr[4323] : arr[4322];
wire r1_2163;
assign r1_2163 = in[0]? arr[4325] : arr[4324];
wire r1_2164;
assign r1_2164 = in[0]? arr[4327] : arr[4326];
wire r1_2165;
assign r1_2165 = in[0]? arr[4329] : arr[4328];
wire r1_2166;
assign r1_2166 = in[0]? arr[4331] : arr[4330];
wire r1_2167;
assign r1_2167 = in[0]? arr[4333] : arr[4332];
wire r1_2168;
assign r1_2168 = in[0]? arr[4335] : arr[4334];
wire r1_2169;
assign r1_2169 = in[0]? arr[4337] : arr[4336];
wire r1_2170;
assign r1_2170 = in[0]? arr[4339] : arr[4338];
wire r1_2171;
assign r1_2171 = in[0]? arr[4341] : arr[4340];
wire r1_2172;
assign r1_2172 = in[0]? arr[4343] : arr[4342];
wire r1_2173;
assign r1_2173 = in[0]? arr[4345] : arr[4344];
wire r1_2174;
assign r1_2174 = in[0]? arr[4347] : arr[4346];
wire r1_2175;
assign r1_2175 = in[0]? arr[4349] : arr[4348];
wire r1_2176;
assign r1_2176 = in[0]? arr[4351] : arr[4350];
wire r1_2177;
assign r1_2177 = in[0]? arr[4353] : arr[4352];
wire r1_2178;
assign r1_2178 = in[0]? arr[4355] : arr[4354];
wire r1_2179;
assign r1_2179 = in[0]? arr[4357] : arr[4356];
wire r1_2180;
assign r1_2180 = in[0]? arr[4359] : arr[4358];
wire r1_2181;
assign r1_2181 = in[0]? arr[4361] : arr[4360];
wire r1_2182;
assign r1_2182 = in[0]? arr[4363] : arr[4362];
wire r1_2183;
assign r1_2183 = in[0]? arr[4365] : arr[4364];
wire r1_2184;
assign r1_2184 = in[0]? arr[4367] : arr[4366];
wire r1_2185;
assign r1_2185 = in[0]? arr[4369] : arr[4368];
wire r1_2186;
assign r1_2186 = in[0]? arr[4371] : arr[4370];
wire r1_2187;
assign r1_2187 = in[0]? arr[4373] : arr[4372];
wire r1_2188;
assign r1_2188 = in[0]? arr[4375] : arr[4374];
wire r1_2189;
assign r1_2189 = in[0]? arr[4377] : arr[4376];
wire r1_2190;
assign r1_2190 = in[0]? arr[4379] : arr[4378];
wire r1_2191;
assign r1_2191 = in[0]? arr[4381] : arr[4380];
wire r1_2192;
assign r1_2192 = in[0]? arr[4383] : arr[4382];
wire r1_2193;
assign r1_2193 = in[0]? arr[4385] : arr[4384];
wire r1_2194;
assign r1_2194 = in[0]? arr[4387] : arr[4386];
wire r1_2195;
assign r1_2195 = in[0]? arr[4389] : arr[4388];
wire r1_2196;
assign r1_2196 = in[0]? arr[4391] : arr[4390];
wire r1_2197;
assign r1_2197 = in[0]? arr[4393] : arr[4392];
wire r1_2198;
assign r1_2198 = in[0]? arr[4395] : arr[4394];
wire r1_2199;
assign r1_2199 = in[0]? arr[4397] : arr[4396];
wire r1_2200;
assign r1_2200 = in[0]? arr[4399] : arr[4398];
wire r1_2201;
assign r1_2201 = in[0]? arr[4401] : arr[4400];
wire r1_2202;
assign r1_2202 = in[0]? arr[4403] : arr[4402];
wire r1_2203;
assign r1_2203 = in[0]? arr[4405] : arr[4404];
wire r1_2204;
assign r1_2204 = in[0]? arr[4407] : arr[4406];
wire r1_2205;
assign r1_2205 = in[0]? arr[4409] : arr[4408];
wire r1_2206;
assign r1_2206 = in[0]? arr[4411] : arr[4410];
wire r1_2207;
assign r1_2207 = in[0]? arr[4413] : arr[4412];
wire r1_2208;
assign r1_2208 = in[0]? arr[4415] : arr[4414];
wire r1_2209;
assign r1_2209 = in[0]? arr[4417] : arr[4416];
wire r1_2210;
assign r1_2210 = in[0]? arr[4419] : arr[4418];
wire r1_2211;
assign r1_2211 = in[0]? arr[4421] : arr[4420];
wire r1_2212;
assign r1_2212 = in[0]? arr[4423] : arr[4422];
wire r1_2213;
assign r1_2213 = in[0]? arr[4425] : arr[4424];
wire r1_2214;
assign r1_2214 = in[0]? arr[4427] : arr[4426];
wire r1_2215;
assign r1_2215 = in[0]? arr[4429] : arr[4428];
wire r1_2216;
assign r1_2216 = in[0]? arr[4431] : arr[4430];
wire r1_2217;
assign r1_2217 = in[0]? arr[4433] : arr[4432];
wire r1_2218;
assign r1_2218 = in[0]? arr[4435] : arr[4434];
wire r1_2219;
assign r1_2219 = in[0]? arr[4437] : arr[4436];
wire r1_2220;
assign r1_2220 = in[0]? arr[4439] : arr[4438];
wire r1_2221;
assign r1_2221 = in[0]? arr[4441] : arr[4440];
wire r1_2222;
assign r1_2222 = in[0]? arr[4443] : arr[4442];
wire r1_2223;
assign r1_2223 = in[0]? arr[4445] : arr[4444];
wire r1_2224;
assign r1_2224 = in[0]? arr[4447] : arr[4446];
wire r1_2225;
assign r1_2225 = in[0]? arr[4449] : arr[4448];
wire r1_2226;
assign r1_2226 = in[0]? arr[4451] : arr[4450];
wire r1_2227;
assign r1_2227 = in[0]? arr[4453] : arr[4452];
wire r1_2228;
assign r1_2228 = in[0]? arr[4455] : arr[4454];
wire r1_2229;
assign r1_2229 = in[0]? arr[4457] : arr[4456];
wire r1_2230;
assign r1_2230 = in[0]? arr[4459] : arr[4458];
wire r1_2231;
assign r1_2231 = in[0]? arr[4461] : arr[4460];
wire r1_2232;
assign r1_2232 = in[0]? arr[4463] : arr[4462];
wire r1_2233;
assign r1_2233 = in[0]? arr[4465] : arr[4464];
wire r1_2234;
assign r1_2234 = in[0]? arr[4467] : arr[4466];
wire r1_2235;
assign r1_2235 = in[0]? arr[4469] : arr[4468];
wire r1_2236;
assign r1_2236 = in[0]? arr[4471] : arr[4470];
wire r1_2237;
assign r1_2237 = in[0]? arr[4473] : arr[4472];
wire r1_2238;
assign r1_2238 = in[0]? arr[4475] : arr[4474];
wire r1_2239;
assign r1_2239 = in[0]? arr[4477] : arr[4476];
wire r1_2240;
assign r1_2240 = in[0]? arr[4479] : arr[4478];
wire r1_2241;
assign r1_2241 = in[0]? arr[4481] : arr[4480];
wire r1_2242;
assign r1_2242 = in[0]? arr[4483] : arr[4482];
wire r1_2243;
assign r1_2243 = in[0]? arr[4485] : arr[4484];
wire r1_2244;
assign r1_2244 = in[0]? arr[4487] : arr[4486];
wire r1_2245;
assign r1_2245 = in[0]? arr[4489] : arr[4488];
wire r1_2246;
assign r1_2246 = in[0]? arr[4491] : arr[4490];
wire r1_2247;
assign r1_2247 = in[0]? arr[4493] : arr[4492];
wire r1_2248;
assign r1_2248 = in[0]? arr[4495] : arr[4494];
wire r1_2249;
assign r1_2249 = in[0]? arr[4497] : arr[4496];
wire r1_2250;
assign r1_2250 = in[0]? arr[4499] : arr[4498];
wire r1_2251;
assign r1_2251 = in[0]? arr[4501] : arr[4500];
wire r1_2252;
assign r1_2252 = in[0]? arr[4503] : arr[4502];
wire r1_2253;
assign r1_2253 = in[0]? arr[4505] : arr[4504];
wire r1_2254;
assign r1_2254 = in[0]? arr[4507] : arr[4506];
wire r1_2255;
assign r1_2255 = in[0]? arr[4509] : arr[4508];
wire r1_2256;
assign r1_2256 = in[0]? arr[4511] : arr[4510];
wire r1_2257;
assign r1_2257 = in[0]? arr[4513] : arr[4512];
wire r1_2258;
assign r1_2258 = in[0]? arr[4515] : arr[4514];
wire r1_2259;
assign r1_2259 = in[0]? arr[4517] : arr[4516];
wire r1_2260;
assign r1_2260 = in[0]? arr[4519] : arr[4518];
wire r1_2261;
assign r1_2261 = in[0]? arr[4521] : arr[4520];
wire r1_2262;
assign r1_2262 = in[0]? arr[4523] : arr[4522];
wire r1_2263;
assign r1_2263 = in[0]? arr[4525] : arr[4524];
wire r1_2264;
assign r1_2264 = in[0]? arr[4527] : arr[4526];
wire r1_2265;
assign r1_2265 = in[0]? arr[4529] : arr[4528];
wire r1_2266;
assign r1_2266 = in[0]? arr[4531] : arr[4530];
wire r1_2267;
assign r1_2267 = in[0]? arr[4533] : arr[4532];
wire r1_2268;
assign r1_2268 = in[0]? arr[4535] : arr[4534];
wire r1_2269;
assign r1_2269 = in[0]? arr[4537] : arr[4536];
wire r1_2270;
assign r1_2270 = in[0]? arr[4539] : arr[4538];
wire r1_2271;
assign r1_2271 = in[0]? arr[4541] : arr[4540];
wire r1_2272;
assign r1_2272 = in[0]? arr[4543] : arr[4542];
wire r1_2273;
assign r1_2273 = in[0]? arr[4545] : arr[4544];
wire r1_2274;
assign r1_2274 = in[0]? arr[4547] : arr[4546];
wire r1_2275;
assign r1_2275 = in[0]? arr[4549] : arr[4548];
wire r1_2276;
assign r1_2276 = in[0]? arr[4551] : arr[4550];
wire r1_2277;
assign r1_2277 = in[0]? arr[4553] : arr[4552];
wire r1_2278;
assign r1_2278 = in[0]? arr[4555] : arr[4554];
wire r1_2279;
assign r1_2279 = in[0]? arr[4557] : arr[4556];
wire r1_2280;
assign r1_2280 = in[0]? arr[4559] : arr[4558];
wire r1_2281;
assign r1_2281 = in[0]? arr[4561] : arr[4560];
wire r1_2282;
assign r1_2282 = in[0]? arr[4563] : arr[4562];
wire r1_2283;
assign r1_2283 = in[0]? arr[4565] : arr[4564];
wire r1_2284;
assign r1_2284 = in[0]? arr[4567] : arr[4566];
wire r1_2285;
assign r1_2285 = in[0]? arr[4569] : arr[4568];
wire r1_2286;
assign r1_2286 = in[0]? arr[4571] : arr[4570];
wire r1_2287;
assign r1_2287 = in[0]? arr[4573] : arr[4572];
wire r1_2288;
assign r1_2288 = in[0]? arr[4575] : arr[4574];
wire r1_2289;
assign r1_2289 = in[0]? arr[4577] : arr[4576];
wire r1_2290;
assign r1_2290 = in[0]? arr[4579] : arr[4578];
wire r1_2291;
assign r1_2291 = in[0]? arr[4581] : arr[4580];
wire r1_2292;
assign r1_2292 = in[0]? arr[4583] : arr[4582];
wire r1_2293;
assign r1_2293 = in[0]? arr[4585] : arr[4584];
wire r1_2294;
assign r1_2294 = in[0]? arr[4587] : arr[4586];
wire r1_2295;
assign r1_2295 = in[0]? arr[4589] : arr[4588];
wire r1_2296;
assign r1_2296 = in[0]? arr[4591] : arr[4590];
wire r1_2297;
assign r1_2297 = in[0]? arr[4593] : arr[4592];
wire r1_2298;
assign r1_2298 = in[0]? arr[4595] : arr[4594];
wire r1_2299;
assign r1_2299 = in[0]? arr[4597] : arr[4596];
wire r1_2300;
assign r1_2300 = in[0]? arr[4599] : arr[4598];
wire r1_2301;
assign r1_2301 = in[0]? arr[4601] : arr[4600];
wire r1_2302;
assign r1_2302 = in[0]? arr[4603] : arr[4602];
wire r1_2303;
assign r1_2303 = in[0]? arr[4605] : arr[4604];
wire r1_2304;
assign r1_2304 = in[0]? arr[4607] : arr[4606];
wire r1_2305;
assign r1_2305 = in[0]? arr[4609] : arr[4608];
wire r1_2306;
assign r1_2306 = in[0]? arr[4611] : arr[4610];
wire r1_2307;
assign r1_2307 = in[0]? arr[4613] : arr[4612];
wire r1_2308;
assign r1_2308 = in[0]? arr[4615] : arr[4614];
wire r1_2309;
assign r1_2309 = in[0]? arr[4617] : arr[4616];
wire r1_2310;
assign r1_2310 = in[0]? arr[4619] : arr[4618];
wire r1_2311;
assign r1_2311 = in[0]? arr[4621] : arr[4620];
wire r1_2312;
assign r1_2312 = in[0]? arr[4623] : arr[4622];
wire r1_2313;
assign r1_2313 = in[0]? arr[4625] : arr[4624];
wire r1_2314;
assign r1_2314 = in[0]? arr[4627] : arr[4626];
wire r1_2315;
assign r1_2315 = in[0]? arr[4629] : arr[4628];
wire r1_2316;
assign r1_2316 = in[0]? arr[4631] : arr[4630];
wire r1_2317;
assign r1_2317 = in[0]? arr[4633] : arr[4632];
wire r1_2318;
assign r1_2318 = in[0]? arr[4635] : arr[4634];
wire r1_2319;
assign r1_2319 = in[0]? arr[4637] : arr[4636];
wire r1_2320;
assign r1_2320 = in[0]? arr[4639] : arr[4638];
wire r1_2321;
assign r1_2321 = in[0]? arr[4641] : arr[4640];
wire r1_2322;
assign r1_2322 = in[0]? arr[4643] : arr[4642];
wire r1_2323;
assign r1_2323 = in[0]? arr[4645] : arr[4644];
wire r1_2324;
assign r1_2324 = in[0]? arr[4647] : arr[4646];
wire r1_2325;
assign r1_2325 = in[0]? arr[4649] : arr[4648];
wire r1_2326;
assign r1_2326 = in[0]? arr[4651] : arr[4650];
wire r1_2327;
assign r1_2327 = in[0]? arr[4653] : arr[4652];
wire r1_2328;
assign r1_2328 = in[0]? arr[4655] : arr[4654];
wire r1_2329;
assign r1_2329 = in[0]? arr[4657] : arr[4656];
wire r1_2330;
assign r1_2330 = in[0]? arr[4659] : arr[4658];
wire r1_2331;
assign r1_2331 = in[0]? arr[4661] : arr[4660];
wire r1_2332;
assign r1_2332 = in[0]? arr[4663] : arr[4662];
wire r1_2333;
assign r1_2333 = in[0]? arr[4665] : arr[4664];
wire r1_2334;
assign r1_2334 = in[0]? arr[4667] : arr[4666];
wire r1_2335;
assign r1_2335 = in[0]? arr[4669] : arr[4668];
wire r1_2336;
assign r1_2336 = in[0]? arr[4671] : arr[4670];
wire r1_2337;
assign r1_2337 = in[0]? arr[4673] : arr[4672];
wire r1_2338;
assign r1_2338 = in[0]? arr[4675] : arr[4674];
wire r1_2339;
assign r1_2339 = in[0]? arr[4677] : arr[4676];
wire r1_2340;
assign r1_2340 = in[0]? arr[4679] : arr[4678];
wire r1_2341;
assign r1_2341 = in[0]? arr[4681] : arr[4680];
wire r1_2342;
assign r1_2342 = in[0]? arr[4683] : arr[4682];
wire r1_2343;
assign r1_2343 = in[0]? arr[4685] : arr[4684];
wire r1_2344;
assign r1_2344 = in[0]? arr[4687] : arr[4686];
wire r1_2345;
assign r1_2345 = in[0]? arr[4689] : arr[4688];
wire r1_2346;
assign r1_2346 = in[0]? arr[4691] : arr[4690];
wire r1_2347;
assign r1_2347 = in[0]? arr[4693] : arr[4692];
wire r1_2348;
assign r1_2348 = in[0]? arr[4695] : arr[4694];
wire r1_2349;
assign r1_2349 = in[0]? arr[4697] : arr[4696];
wire r1_2350;
assign r1_2350 = in[0]? arr[4699] : arr[4698];
wire r1_2351;
assign r1_2351 = in[0]? arr[4701] : arr[4700];
wire r1_2352;
assign r1_2352 = in[0]? arr[4703] : arr[4702];
wire r1_2353;
assign r1_2353 = in[0]? arr[4705] : arr[4704];
wire r1_2354;
assign r1_2354 = in[0]? arr[4707] : arr[4706];
wire r1_2355;
assign r1_2355 = in[0]? arr[4709] : arr[4708];
wire r1_2356;
assign r1_2356 = in[0]? arr[4711] : arr[4710];
wire r1_2357;
assign r1_2357 = in[0]? arr[4713] : arr[4712];
wire r1_2358;
assign r1_2358 = in[0]? arr[4715] : arr[4714];
wire r1_2359;
assign r1_2359 = in[0]? arr[4717] : arr[4716];
wire r1_2360;
assign r1_2360 = in[0]? arr[4719] : arr[4718];
wire r1_2361;
assign r1_2361 = in[0]? arr[4721] : arr[4720];
wire r1_2362;
assign r1_2362 = in[0]? arr[4723] : arr[4722];
wire r1_2363;
assign r1_2363 = in[0]? arr[4725] : arr[4724];
wire r1_2364;
assign r1_2364 = in[0]? arr[4727] : arr[4726];
wire r1_2365;
assign r1_2365 = in[0]? arr[4729] : arr[4728];
wire r1_2366;
assign r1_2366 = in[0]? arr[4731] : arr[4730];
wire r1_2367;
assign r1_2367 = in[0]? arr[4733] : arr[4732];
wire r1_2368;
assign r1_2368 = in[0]? arr[4735] : arr[4734];
wire r1_2369;
assign r1_2369 = in[0]? arr[4737] : arr[4736];
wire r1_2370;
assign r1_2370 = in[0]? arr[4739] : arr[4738];
wire r1_2371;
assign r1_2371 = in[0]? arr[4741] : arr[4740];
wire r1_2372;
assign r1_2372 = in[0]? arr[4743] : arr[4742];
wire r1_2373;
assign r1_2373 = in[0]? arr[4745] : arr[4744];
wire r1_2374;
assign r1_2374 = in[0]? arr[4747] : arr[4746];
wire r1_2375;
assign r1_2375 = in[0]? arr[4749] : arr[4748];
wire r1_2376;
assign r1_2376 = in[0]? arr[4751] : arr[4750];
wire r1_2377;
assign r1_2377 = in[0]? arr[4753] : arr[4752];
wire r1_2378;
assign r1_2378 = in[0]? arr[4755] : arr[4754];
wire r1_2379;
assign r1_2379 = in[0]? arr[4757] : arr[4756];
wire r1_2380;
assign r1_2380 = in[0]? arr[4759] : arr[4758];
wire r1_2381;
assign r1_2381 = in[0]? arr[4761] : arr[4760];
wire r1_2382;
assign r1_2382 = in[0]? arr[4763] : arr[4762];
wire r1_2383;
assign r1_2383 = in[0]? arr[4765] : arr[4764];
wire r1_2384;
assign r1_2384 = in[0]? arr[4767] : arr[4766];
wire r1_2385;
assign r1_2385 = in[0]? arr[4769] : arr[4768];
wire r1_2386;
assign r1_2386 = in[0]? arr[4771] : arr[4770];
wire r1_2387;
assign r1_2387 = in[0]? arr[4773] : arr[4772];
wire r1_2388;
assign r1_2388 = in[0]? arr[4775] : arr[4774];
wire r1_2389;
assign r1_2389 = in[0]? arr[4777] : arr[4776];
wire r1_2390;
assign r1_2390 = in[0]? arr[4779] : arr[4778];
wire r1_2391;
assign r1_2391 = in[0]? arr[4781] : arr[4780];
wire r1_2392;
assign r1_2392 = in[0]? arr[4783] : arr[4782];
wire r1_2393;
assign r1_2393 = in[0]? arr[4785] : arr[4784];
wire r1_2394;
assign r1_2394 = in[0]? arr[4787] : arr[4786];
wire r1_2395;
assign r1_2395 = in[0]? arr[4789] : arr[4788];
wire r1_2396;
assign r1_2396 = in[0]? arr[4791] : arr[4790];
wire r1_2397;
assign r1_2397 = in[0]? arr[4793] : arr[4792];
wire r1_2398;
assign r1_2398 = in[0]? arr[4795] : arr[4794];
wire r1_2399;
assign r1_2399 = in[0]? arr[4797] : arr[4796];
wire r1_2400;
assign r1_2400 = in[0]? arr[4799] : arr[4798];
wire r1_2401;
assign r1_2401 = in[0]? arr[4801] : arr[4800];
wire r1_2402;
assign r1_2402 = in[0]? arr[4803] : arr[4802];
wire r1_2403;
assign r1_2403 = in[0]? arr[4805] : arr[4804];
wire r1_2404;
assign r1_2404 = in[0]? arr[4807] : arr[4806];
wire r1_2405;
assign r1_2405 = in[0]? arr[4809] : arr[4808];
wire r1_2406;
assign r1_2406 = in[0]? arr[4811] : arr[4810];
wire r1_2407;
assign r1_2407 = in[0]? arr[4813] : arr[4812];
wire r1_2408;
assign r1_2408 = in[0]? arr[4815] : arr[4814];
wire r1_2409;
assign r1_2409 = in[0]? arr[4817] : arr[4816];
wire r1_2410;
assign r1_2410 = in[0]? arr[4819] : arr[4818];
wire r1_2411;
assign r1_2411 = in[0]? arr[4821] : arr[4820];
wire r1_2412;
assign r1_2412 = in[0]? arr[4823] : arr[4822];
wire r1_2413;
assign r1_2413 = in[0]? arr[4825] : arr[4824];
wire r1_2414;
assign r1_2414 = in[0]? arr[4827] : arr[4826];
wire r1_2415;
assign r1_2415 = in[0]? arr[4829] : arr[4828];
wire r1_2416;
assign r1_2416 = in[0]? arr[4831] : arr[4830];
wire r1_2417;
assign r1_2417 = in[0]? arr[4833] : arr[4832];
wire r1_2418;
assign r1_2418 = in[0]? arr[4835] : arr[4834];
wire r1_2419;
assign r1_2419 = in[0]? arr[4837] : arr[4836];
wire r1_2420;
assign r1_2420 = in[0]? arr[4839] : arr[4838];
wire r1_2421;
assign r1_2421 = in[0]? arr[4841] : arr[4840];
wire r1_2422;
assign r1_2422 = in[0]? arr[4843] : arr[4842];
wire r1_2423;
assign r1_2423 = in[0]? arr[4845] : arr[4844];
wire r1_2424;
assign r1_2424 = in[0]? arr[4847] : arr[4846];
wire r1_2425;
assign r1_2425 = in[0]? arr[4849] : arr[4848];
wire r1_2426;
assign r1_2426 = in[0]? arr[4851] : arr[4850];
wire r1_2427;
assign r1_2427 = in[0]? arr[4853] : arr[4852];
wire r1_2428;
assign r1_2428 = in[0]? arr[4855] : arr[4854];
wire r1_2429;
assign r1_2429 = in[0]? arr[4857] : arr[4856];
wire r1_2430;
assign r1_2430 = in[0]? arr[4859] : arr[4858];
wire r1_2431;
assign r1_2431 = in[0]? arr[4861] : arr[4860];
wire r1_2432;
assign r1_2432 = in[0]? arr[4863] : arr[4862];
wire r1_2433;
assign r1_2433 = in[0]? arr[4865] : arr[4864];
wire r1_2434;
assign r1_2434 = in[0]? arr[4867] : arr[4866];
wire r1_2435;
assign r1_2435 = in[0]? arr[4869] : arr[4868];
wire r1_2436;
assign r1_2436 = in[0]? arr[4871] : arr[4870];
wire r1_2437;
assign r1_2437 = in[0]? arr[4873] : arr[4872];
wire r1_2438;
assign r1_2438 = in[0]? arr[4875] : arr[4874];
wire r1_2439;
assign r1_2439 = in[0]? arr[4877] : arr[4876];
wire r1_2440;
assign r1_2440 = in[0]? arr[4879] : arr[4878];
wire r1_2441;
assign r1_2441 = in[0]? arr[4881] : arr[4880];
wire r1_2442;
assign r1_2442 = in[0]? arr[4883] : arr[4882];
wire r1_2443;
assign r1_2443 = in[0]? arr[4885] : arr[4884];
wire r1_2444;
assign r1_2444 = in[0]? arr[4887] : arr[4886];
wire r1_2445;
assign r1_2445 = in[0]? arr[4889] : arr[4888];
wire r1_2446;
assign r1_2446 = in[0]? arr[4891] : arr[4890];
wire r1_2447;
assign r1_2447 = in[0]? arr[4893] : arr[4892];
wire r1_2448;
assign r1_2448 = in[0]? arr[4895] : arr[4894];
wire r1_2449;
assign r1_2449 = in[0]? arr[4897] : arr[4896];
wire r1_2450;
assign r1_2450 = in[0]? arr[4899] : arr[4898];
wire r1_2451;
assign r1_2451 = in[0]? arr[4901] : arr[4900];
wire r1_2452;
assign r1_2452 = in[0]? arr[4903] : arr[4902];
wire r1_2453;
assign r1_2453 = in[0]? arr[4905] : arr[4904];
wire r1_2454;
assign r1_2454 = in[0]? arr[4907] : arr[4906];
wire r1_2455;
assign r1_2455 = in[0]? arr[4909] : arr[4908];
wire r1_2456;
assign r1_2456 = in[0]? arr[4911] : arr[4910];
wire r1_2457;
assign r1_2457 = in[0]? arr[4913] : arr[4912];
wire r1_2458;
assign r1_2458 = in[0]? arr[4915] : arr[4914];
wire r1_2459;
assign r1_2459 = in[0]? arr[4917] : arr[4916];
wire r1_2460;
assign r1_2460 = in[0]? arr[4919] : arr[4918];
wire r1_2461;
assign r1_2461 = in[0]? arr[4921] : arr[4920];
wire r1_2462;
assign r1_2462 = in[0]? arr[4923] : arr[4922];
wire r1_2463;
assign r1_2463 = in[0]? arr[4925] : arr[4924];
wire r1_2464;
assign r1_2464 = in[0]? arr[4927] : arr[4926];
wire r1_2465;
assign r1_2465 = in[0]? arr[4929] : arr[4928];
wire r1_2466;
assign r1_2466 = in[0]? arr[4931] : arr[4930];
wire r1_2467;
assign r1_2467 = in[0]? arr[4933] : arr[4932];
wire r1_2468;
assign r1_2468 = in[0]? arr[4935] : arr[4934];
wire r1_2469;
assign r1_2469 = in[0]? arr[4937] : arr[4936];
wire r1_2470;
assign r1_2470 = in[0]? arr[4939] : arr[4938];
wire r1_2471;
assign r1_2471 = in[0]? arr[4941] : arr[4940];
wire r1_2472;
assign r1_2472 = in[0]? arr[4943] : arr[4942];
wire r1_2473;
assign r1_2473 = in[0]? arr[4945] : arr[4944];
wire r1_2474;
assign r1_2474 = in[0]? arr[4947] : arr[4946];
wire r1_2475;
assign r1_2475 = in[0]? arr[4949] : arr[4948];
wire r1_2476;
assign r1_2476 = in[0]? arr[4951] : arr[4950];
wire r1_2477;
assign r1_2477 = in[0]? arr[4953] : arr[4952];
wire r1_2478;
assign r1_2478 = in[0]? arr[4955] : arr[4954];
wire r1_2479;
assign r1_2479 = in[0]? arr[4957] : arr[4956];
wire r1_2480;
assign r1_2480 = in[0]? arr[4959] : arr[4958];
wire r1_2481;
assign r1_2481 = in[0]? arr[4961] : arr[4960];
wire r1_2482;
assign r1_2482 = in[0]? arr[4963] : arr[4962];
wire r1_2483;
assign r1_2483 = in[0]? arr[4965] : arr[4964];
wire r1_2484;
assign r1_2484 = in[0]? arr[4967] : arr[4966];
wire r1_2485;
assign r1_2485 = in[0]? arr[4969] : arr[4968];
wire r1_2486;
assign r1_2486 = in[0]? arr[4971] : arr[4970];
wire r1_2487;
assign r1_2487 = in[0]? arr[4973] : arr[4972];
wire r1_2488;
assign r1_2488 = in[0]? arr[4975] : arr[4974];
wire r1_2489;
assign r1_2489 = in[0]? arr[4977] : arr[4976];
wire r1_2490;
assign r1_2490 = in[0]? arr[4979] : arr[4978];
wire r1_2491;
assign r1_2491 = in[0]? arr[4981] : arr[4980];
wire r1_2492;
assign r1_2492 = in[0]? arr[4983] : arr[4982];
wire r1_2493;
assign r1_2493 = in[0]? arr[4985] : arr[4984];
wire r1_2494;
assign r1_2494 = in[0]? arr[4987] : arr[4986];
wire r1_2495;
assign r1_2495 = in[0]? arr[4989] : arr[4988];
wire r1_2496;
assign r1_2496 = in[0]? arr[4991] : arr[4990];
wire r1_2497;
assign r1_2497 = in[0]? arr[4993] : arr[4992];
wire r1_2498;
assign r1_2498 = in[0]? arr[4995] : arr[4994];
wire r1_2499;
assign r1_2499 = in[0]? arr[4997] : arr[4996];
wire r1_2500;
assign r1_2500 = in[0]? arr[4999] : arr[4998];
wire r1_2501;
assign r1_2501 = in[0]? arr[5001] : arr[5000];
wire r1_2502;
assign r1_2502 = in[0]? arr[5003] : arr[5002];
wire r1_2503;
assign r1_2503 = in[0]? arr[5005] : arr[5004];
wire r1_2504;
assign r1_2504 = in[0]? arr[5007] : arr[5006];
wire r1_2505;
assign r1_2505 = in[0]? arr[5009] : arr[5008];
wire r1_2506;
assign r1_2506 = in[0]? arr[5011] : arr[5010];
wire r1_2507;
assign r1_2507 = in[0]? arr[5013] : arr[5012];
wire r1_2508;
assign r1_2508 = in[0]? arr[5015] : arr[5014];
wire r1_2509;
assign r1_2509 = in[0]? arr[5017] : arr[5016];
wire r1_2510;
assign r1_2510 = in[0]? arr[5019] : arr[5018];
wire r1_2511;
assign r1_2511 = in[0]? arr[5021] : arr[5020];
wire r1_2512;
assign r1_2512 = in[0]? arr[5023] : arr[5022];
wire r1_2513;
assign r1_2513 = in[0]? arr[5025] : arr[5024];
wire r1_2514;
assign r1_2514 = in[0]? arr[5027] : arr[5026];
wire r1_2515;
assign r1_2515 = in[0]? arr[5029] : arr[5028];
wire r1_2516;
assign r1_2516 = in[0]? arr[5031] : arr[5030];
wire r1_2517;
assign r1_2517 = in[0]? arr[5033] : arr[5032];
wire r1_2518;
assign r1_2518 = in[0]? arr[5035] : arr[5034];
wire r1_2519;
assign r1_2519 = in[0]? arr[5037] : arr[5036];
wire r1_2520;
assign r1_2520 = in[0]? arr[5039] : arr[5038];
wire r1_2521;
assign r1_2521 = in[0]? arr[5041] : arr[5040];
wire r1_2522;
assign r1_2522 = in[0]? arr[5043] : arr[5042];
wire r1_2523;
assign r1_2523 = in[0]? arr[5045] : arr[5044];
wire r1_2524;
assign r1_2524 = in[0]? arr[5047] : arr[5046];
wire r1_2525;
assign r1_2525 = in[0]? arr[5049] : arr[5048];
wire r1_2526;
assign r1_2526 = in[0]? arr[5051] : arr[5050];
wire r1_2527;
assign r1_2527 = in[0]? arr[5053] : arr[5052];
wire r1_2528;
assign r1_2528 = in[0]? arr[5055] : arr[5054];
wire r1_2529;
assign r1_2529 = in[0]? arr[5057] : arr[5056];
wire r1_2530;
assign r1_2530 = in[0]? arr[5059] : arr[5058];
wire r1_2531;
assign r1_2531 = in[0]? arr[5061] : arr[5060];
wire r1_2532;
assign r1_2532 = in[0]? arr[5063] : arr[5062];
wire r1_2533;
assign r1_2533 = in[0]? arr[5065] : arr[5064];
wire r1_2534;
assign r1_2534 = in[0]? arr[5067] : arr[5066];
wire r1_2535;
assign r1_2535 = in[0]? arr[5069] : arr[5068];
wire r1_2536;
assign r1_2536 = in[0]? arr[5071] : arr[5070];
wire r1_2537;
assign r1_2537 = in[0]? arr[5073] : arr[5072];
wire r1_2538;
assign r1_2538 = in[0]? arr[5075] : arr[5074];
wire r1_2539;
assign r1_2539 = in[0]? arr[5077] : arr[5076];
wire r1_2540;
assign r1_2540 = in[0]? arr[5079] : arr[5078];
wire r1_2541;
assign r1_2541 = in[0]? arr[5081] : arr[5080];
wire r1_2542;
assign r1_2542 = in[0]? arr[5083] : arr[5082];
wire r1_2543;
assign r1_2543 = in[0]? arr[5085] : arr[5084];
wire r1_2544;
assign r1_2544 = in[0]? arr[5087] : arr[5086];
wire r1_2545;
assign r1_2545 = in[0]? arr[5089] : arr[5088];
wire r1_2546;
assign r1_2546 = in[0]? arr[5091] : arr[5090];
wire r1_2547;
assign r1_2547 = in[0]? arr[5093] : arr[5092];
wire r1_2548;
assign r1_2548 = in[0]? arr[5095] : arr[5094];
wire r1_2549;
assign r1_2549 = in[0]? arr[5097] : arr[5096];
wire r1_2550;
assign r1_2550 = in[0]? arr[5099] : arr[5098];
wire r1_2551;
assign r1_2551 = in[0]? arr[5101] : arr[5100];
wire r1_2552;
assign r1_2552 = in[0]? arr[5103] : arr[5102];
wire r1_2553;
assign r1_2553 = in[0]? arr[5105] : arr[5104];
wire r1_2554;
assign r1_2554 = in[0]? arr[5107] : arr[5106];
wire r1_2555;
assign r1_2555 = in[0]? arr[5109] : arr[5108];
wire r1_2556;
assign r1_2556 = in[0]? arr[5111] : arr[5110];
wire r1_2557;
assign r1_2557 = in[0]? arr[5113] : arr[5112];
wire r1_2558;
assign r1_2558 = in[0]? arr[5115] : arr[5114];
wire r1_2559;
assign r1_2559 = in[0]? arr[5117] : arr[5116];
wire r1_2560;
assign r1_2560 = in[0]? arr[5119] : arr[5118];
wire r1_2561;
assign r1_2561 = in[0]? arr[5121] : arr[5120];
wire r1_2562;
assign r1_2562 = in[0]? arr[5123] : arr[5122];
wire r1_2563;
assign r1_2563 = in[0]? arr[5125] : arr[5124];
wire r1_2564;
assign r1_2564 = in[0]? arr[5127] : arr[5126];
wire r1_2565;
assign r1_2565 = in[0]? arr[5129] : arr[5128];
wire r1_2566;
assign r1_2566 = in[0]? arr[5131] : arr[5130];
wire r1_2567;
assign r1_2567 = in[0]? arr[5133] : arr[5132];
wire r1_2568;
assign r1_2568 = in[0]? arr[5135] : arr[5134];
wire r1_2569;
assign r1_2569 = in[0]? arr[5137] : arr[5136];
wire r1_2570;
assign r1_2570 = in[0]? arr[5139] : arr[5138];
wire r1_2571;
assign r1_2571 = in[0]? arr[5141] : arr[5140];
wire r1_2572;
assign r1_2572 = in[0]? arr[5143] : arr[5142];
wire r1_2573;
assign r1_2573 = in[0]? arr[5145] : arr[5144];
wire r1_2574;
assign r1_2574 = in[0]? arr[5147] : arr[5146];
wire r1_2575;
assign r1_2575 = in[0]? arr[5149] : arr[5148];
wire r1_2576;
assign r1_2576 = in[0]? arr[5151] : arr[5150];
wire r1_2577;
assign r1_2577 = in[0]? arr[5153] : arr[5152];
wire r1_2578;
assign r1_2578 = in[0]? arr[5155] : arr[5154];
wire r1_2579;
assign r1_2579 = in[0]? arr[5157] : arr[5156];
wire r1_2580;
assign r1_2580 = in[0]? arr[5159] : arr[5158];
wire r1_2581;
assign r1_2581 = in[0]? arr[5161] : arr[5160];
wire r1_2582;
assign r1_2582 = in[0]? arr[5163] : arr[5162];
wire r1_2583;
assign r1_2583 = in[0]? arr[5165] : arr[5164];
wire r1_2584;
assign r1_2584 = in[0]? arr[5167] : arr[5166];
wire r1_2585;
assign r1_2585 = in[0]? arr[5169] : arr[5168];
wire r1_2586;
assign r1_2586 = in[0]? arr[5171] : arr[5170];
wire r1_2587;
assign r1_2587 = in[0]? arr[5173] : arr[5172];
wire r1_2588;
assign r1_2588 = in[0]? arr[5175] : arr[5174];
wire r1_2589;
assign r1_2589 = in[0]? arr[5177] : arr[5176];
wire r1_2590;
assign r1_2590 = in[0]? arr[5179] : arr[5178];
wire r1_2591;
assign r1_2591 = in[0]? arr[5181] : arr[5180];
wire r1_2592;
assign r1_2592 = in[0]? arr[5183] : arr[5182];
wire r1_2593;
assign r1_2593 = in[0]? arr[5185] : arr[5184];
wire r1_2594;
assign r1_2594 = in[0]? arr[5187] : arr[5186];
wire r1_2595;
assign r1_2595 = in[0]? arr[5189] : arr[5188];
wire r1_2596;
assign r1_2596 = in[0]? arr[5191] : arr[5190];
wire r1_2597;
assign r1_2597 = in[0]? arr[5193] : arr[5192];
wire r1_2598;
assign r1_2598 = in[0]? arr[5195] : arr[5194];
wire r1_2599;
assign r1_2599 = in[0]? arr[5197] : arr[5196];
wire r1_2600;
assign r1_2600 = in[0]? arr[5199] : arr[5198];
wire r1_2601;
assign r1_2601 = in[0]? arr[5201] : arr[5200];
wire r1_2602;
assign r1_2602 = in[0]? arr[5203] : arr[5202];
wire r1_2603;
assign r1_2603 = in[0]? arr[5205] : arr[5204];
wire r1_2604;
assign r1_2604 = in[0]? arr[5207] : arr[5206];
wire r1_2605;
assign r1_2605 = in[0]? arr[5209] : arr[5208];
wire r1_2606;
assign r1_2606 = in[0]? arr[5211] : arr[5210];
wire r1_2607;
assign r1_2607 = in[0]? arr[5213] : arr[5212];
wire r1_2608;
assign r1_2608 = in[0]? arr[5215] : arr[5214];
wire r1_2609;
assign r1_2609 = in[0]? arr[5217] : arr[5216];
wire r1_2610;
assign r1_2610 = in[0]? arr[5219] : arr[5218];
wire r1_2611;
assign r1_2611 = in[0]? arr[5221] : arr[5220];
wire r1_2612;
assign r1_2612 = in[0]? arr[5223] : arr[5222];
wire r1_2613;
assign r1_2613 = in[0]? arr[5225] : arr[5224];
wire r1_2614;
assign r1_2614 = in[0]? arr[5227] : arr[5226];
wire r1_2615;
assign r1_2615 = in[0]? arr[5229] : arr[5228];
wire r1_2616;
assign r1_2616 = in[0]? arr[5231] : arr[5230];
wire r1_2617;
assign r1_2617 = in[0]? arr[5233] : arr[5232];
wire r1_2618;
assign r1_2618 = in[0]? arr[5235] : arr[5234];
wire r1_2619;
assign r1_2619 = in[0]? arr[5237] : arr[5236];
wire r1_2620;
assign r1_2620 = in[0]? arr[5239] : arr[5238];
wire r1_2621;
assign r1_2621 = in[0]? arr[5241] : arr[5240];
wire r1_2622;
assign r1_2622 = in[0]? arr[5243] : arr[5242];
wire r1_2623;
assign r1_2623 = in[0]? arr[5245] : arr[5244];
wire r1_2624;
assign r1_2624 = in[0]? arr[5247] : arr[5246];
wire r1_2625;
assign r1_2625 = in[0]? arr[5249] : arr[5248];
wire r1_2626;
assign r1_2626 = in[0]? arr[5251] : arr[5250];
wire r1_2627;
assign r1_2627 = in[0]? arr[5253] : arr[5252];
wire r1_2628;
assign r1_2628 = in[0]? arr[5255] : arr[5254];
wire r1_2629;
assign r1_2629 = in[0]? arr[5257] : arr[5256];
wire r1_2630;
assign r1_2630 = in[0]? arr[5259] : arr[5258];
wire r1_2631;
assign r1_2631 = in[0]? arr[5261] : arr[5260];
wire r1_2632;
assign r1_2632 = in[0]? arr[5263] : arr[5262];
wire r1_2633;
assign r1_2633 = in[0]? arr[5265] : arr[5264];
wire r1_2634;
assign r1_2634 = in[0]? arr[5267] : arr[5266];
wire r1_2635;
assign r1_2635 = in[0]? arr[5269] : arr[5268];
wire r1_2636;
assign r1_2636 = in[0]? arr[5271] : arr[5270];
wire r1_2637;
assign r1_2637 = in[0]? arr[5273] : arr[5272];
wire r1_2638;
assign r1_2638 = in[0]? arr[5275] : arr[5274];
wire r1_2639;
assign r1_2639 = in[0]? arr[5277] : arr[5276];
wire r1_2640;
assign r1_2640 = in[0]? arr[5279] : arr[5278];
wire r1_2641;
assign r1_2641 = in[0]? arr[5281] : arr[5280];
wire r1_2642;
assign r1_2642 = in[0]? arr[5283] : arr[5282];
wire r1_2643;
assign r1_2643 = in[0]? arr[5285] : arr[5284];
wire r1_2644;
assign r1_2644 = in[0]? arr[5287] : arr[5286];
wire r1_2645;
assign r1_2645 = in[0]? arr[5289] : arr[5288];
wire r1_2646;
assign r1_2646 = in[0]? arr[5291] : arr[5290];
wire r1_2647;
assign r1_2647 = in[0]? arr[5293] : arr[5292];
wire r1_2648;
assign r1_2648 = in[0]? arr[5295] : arr[5294];
wire r1_2649;
assign r1_2649 = in[0]? arr[5297] : arr[5296];
wire r1_2650;
assign r1_2650 = in[0]? arr[5299] : arr[5298];
wire r1_2651;
assign r1_2651 = in[0]? arr[5301] : arr[5300];
wire r1_2652;
assign r1_2652 = in[0]? arr[5303] : arr[5302];
wire r1_2653;
assign r1_2653 = in[0]? arr[5305] : arr[5304];
wire r1_2654;
assign r1_2654 = in[0]? arr[5307] : arr[5306];
wire r1_2655;
assign r1_2655 = in[0]? arr[5309] : arr[5308];
wire r1_2656;
assign r1_2656 = in[0]? arr[5311] : arr[5310];
wire r1_2657;
assign r1_2657 = in[0]? arr[5313] : arr[5312];
wire r1_2658;
assign r1_2658 = in[0]? arr[5315] : arr[5314];
wire r1_2659;
assign r1_2659 = in[0]? arr[5317] : arr[5316];
wire r1_2660;
assign r1_2660 = in[0]? arr[5319] : arr[5318];
wire r1_2661;
assign r1_2661 = in[0]? arr[5321] : arr[5320];
wire r1_2662;
assign r1_2662 = in[0]? arr[5323] : arr[5322];
wire r1_2663;
assign r1_2663 = in[0]? arr[5325] : arr[5324];
wire r1_2664;
assign r1_2664 = in[0]? arr[5327] : arr[5326];
wire r1_2665;
assign r1_2665 = in[0]? arr[5329] : arr[5328];
wire r1_2666;
assign r1_2666 = in[0]? arr[5331] : arr[5330];
wire r1_2667;
assign r1_2667 = in[0]? arr[5333] : arr[5332];
wire r1_2668;
assign r1_2668 = in[0]? arr[5335] : arr[5334];
wire r1_2669;
assign r1_2669 = in[0]? arr[5337] : arr[5336];
wire r1_2670;
assign r1_2670 = in[0]? arr[5339] : arr[5338];
wire r1_2671;
assign r1_2671 = in[0]? arr[5341] : arr[5340];
wire r1_2672;
assign r1_2672 = in[0]? arr[5343] : arr[5342];
wire r1_2673;
assign r1_2673 = in[0]? arr[5345] : arr[5344];
wire r1_2674;
assign r1_2674 = in[0]? arr[5347] : arr[5346];
wire r1_2675;
assign r1_2675 = in[0]? arr[5349] : arr[5348];
wire r1_2676;
assign r1_2676 = in[0]? arr[5351] : arr[5350];
wire r1_2677;
assign r1_2677 = in[0]? arr[5353] : arr[5352];
wire r1_2678;
assign r1_2678 = in[0]? arr[5355] : arr[5354];
wire r1_2679;
assign r1_2679 = in[0]? arr[5357] : arr[5356];
wire r1_2680;
assign r1_2680 = in[0]? arr[5359] : arr[5358];
wire r1_2681;
assign r1_2681 = in[0]? arr[5361] : arr[5360];
wire r1_2682;
assign r1_2682 = in[0]? arr[5363] : arr[5362];
wire r1_2683;
assign r1_2683 = in[0]? arr[5365] : arr[5364];
wire r1_2684;
assign r1_2684 = in[0]? arr[5367] : arr[5366];
wire r1_2685;
assign r1_2685 = in[0]? arr[5369] : arr[5368];
wire r1_2686;
assign r1_2686 = in[0]? arr[5371] : arr[5370];
wire r1_2687;
assign r1_2687 = in[0]? arr[5373] : arr[5372];
wire r1_2688;
assign r1_2688 = in[0]? arr[5375] : arr[5374];
wire r1_2689;
assign r1_2689 = in[0]? arr[5377] : arr[5376];
wire r1_2690;
assign r1_2690 = in[0]? arr[5379] : arr[5378];
wire r1_2691;
assign r1_2691 = in[0]? arr[5381] : arr[5380];
wire r1_2692;
assign r1_2692 = in[0]? arr[5383] : arr[5382];
wire r1_2693;
assign r1_2693 = in[0]? arr[5385] : arr[5384];
wire r1_2694;
assign r1_2694 = in[0]? arr[5387] : arr[5386];
wire r1_2695;
assign r1_2695 = in[0]? arr[5389] : arr[5388];
wire r1_2696;
assign r1_2696 = in[0]? arr[5391] : arr[5390];
wire r1_2697;
assign r1_2697 = in[0]? arr[5393] : arr[5392];
wire r1_2698;
assign r1_2698 = in[0]? arr[5395] : arr[5394];
wire r1_2699;
assign r1_2699 = in[0]? arr[5397] : arr[5396];
wire r1_2700;
assign r1_2700 = in[0]? arr[5399] : arr[5398];
wire r1_2701;
assign r1_2701 = in[0]? arr[5401] : arr[5400];
wire r1_2702;
assign r1_2702 = in[0]? arr[5403] : arr[5402];
wire r1_2703;
assign r1_2703 = in[0]? arr[5405] : arr[5404];
wire r1_2704;
assign r1_2704 = in[0]? arr[5407] : arr[5406];
wire r1_2705;
assign r1_2705 = in[0]? arr[5409] : arr[5408];
wire r1_2706;
assign r1_2706 = in[0]? arr[5411] : arr[5410];
wire r1_2707;
assign r1_2707 = in[0]? arr[5413] : arr[5412];
wire r1_2708;
assign r1_2708 = in[0]? arr[5415] : arr[5414];
wire r1_2709;
assign r1_2709 = in[0]? arr[5417] : arr[5416];
wire r1_2710;
assign r1_2710 = in[0]? arr[5419] : arr[5418];
wire r1_2711;
assign r1_2711 = in[0]? arr[5421] : arr[5420];
wire r1_2712;
assign r1_2712 = in[0]? arr[5423] : arr[5422];
wire r1_2713;
assign r1_2713 = in[0]? arr[5425] : arr[5424];
wire r1_2714;
assign r1_2714 = in[0]? arr[5427] : arr[5426];
wire r1_2715;
assign r1_2715 = in[0]? arr[5429] : arr[5428];
wire r1_2716;
assign r1_2716 = in[0]? arr[5431] : arr[5430];
wire r1_2717;
assign r1_2717 = in[0]? arr[5433] : arr[5432];
wire r1_2718;
assign r1_2718 = in[0]? arr[5435] : arr[5434];
wire r1_2719;
assign r1_2719 = in[0]? arr[5437] : arr[5436];
wire r1_2720;
assign r1_2720 = in[0]? arr[5439] : arr[5438];
wire r1_2721;
assign r1_2721 = in[0]? arr[5441] : arr[5440];
wire r1_2722;
assign r1_2722 = in[0]? arr[5443] : arr[5442];
wire r1_2723;
assign r1_2723 = in[0]? arr[5445] : arr[5444];
wire r1_2724;
assign r1_2724 = in[0]? arr[5447] : arr[5446];
wire r1_2725;
assign r1_2725 = in[0]? arr[5449] : arr[5448];
wire r1_2726;
assign r1_2726 = in[0]? arr[5451] : arr[5450];
wire r1_2727;
assign r1_2727 = in[0]? arr[5453] : arr[5452];
wire r1_2728;
assign r1_2728 = in[0]? arr[5455] : arr[5454];
wire r1_2729;
assign r1_2729 = in[0]? arr[5457] : arr[5456];
wire r1_2730;
assign r1_2730 = in[0]? arr[5459] : arr[5458];
wire r1_2731;
assign r1_2731 = in[0]? arr[5461] : arr[5460];
wire r1_2732;
assign r1_2732 = in[0]? arr[5463] : arr[5462];
wire r1_2733;
assign r1_2733 = in[0]? arr[5465] : arr[5464];
wire r1_2734;
assign r1_2734 = in[0]? arr[5467] : arr[5466];
wire r1_2735;
assign r1_2735 = in[0]? arr[5469] : arr[5468];
wire r1_2736;
assign r1_2736 = in[0]? arr[5471] : arr[5470];
wire r1_2737;
assign r1_2737 = in[0]? arr[5473] : arr[5472];
wire r1_2738;
assign r1_2738 = in[0]? arr[5475] : arr[5474];
wire r1_2739;
assign r1_2739 = in[0]? arr[5477] : arr[5476];
wire r1_2740;
assign r1_2740 = in[0]? arr[5479] : arr[5478];
wire r1_2741;
assign r1_2741 = in[0]? arr[5481] : arr[5480];
wire r1_2742;
assign r1_2742 = in[0]? arr[5483] : arr[5482];
wire r1_2743;
assign r1_2743 = in[0]? arr[5485] : arr[5484];
wire r1_2744;
assign r1_2744 = in[0]? arr[5487] : arr[5486];
wire r1_2745;
assign r1_2745 = in[0]? arr[5489] : arr[5488];
wire r1_2746;
assign r1_2746 = in[0]? arr[5491] : arr[5490];
wire r1_2747;
assign r1_2747 = in[0]? arr[5493] : arr[5492];
wire r1_2748;
assign r1_2748 = in[0]? arr[5495] : arr[5494];
wire r1_2749;
assign r1_2749 = in[0]? arr[5497] : arr[5496];
wire r1_2750;
assign r1_2750 = in[0]? arr[5499] : arr[5498];
wire r1_2751;
assign r1_2751 = in[0]? arr[5501] : arr[5500];
wire r1_2752;
assign r1_2752 = in[0]? arr[5503] : arr[5502];
wire r1_2753;
assign r1_2753 = in[0]? arr[5505] : arr[5504];
wire r1_2754;
assign r1_2754 = in[0]? arr[5507] : arr[5506];
wire r1_2755;
assign r1_2755 = in[0]? arr[5509] : arr[5508];
wire r1_2756;
assign r1_2756 = in[0]? arr[5511] : arr[5510];
wire r1_2757;
assign r1_2757 = in[0]? arr[5513] : arr[5512];
wire r1_2758;
assign r1_2758 = in[0]? arr[5515] : arr[5514];
wire r1_2759;
assign r1_2759 = in[0]? arr[5517] : arr[5516];
wire r1_2760;
assign r1_2760 = in[0]? arr[5519] : arr[5518];
wire r1_2761;
assign r1_2761 = in[0]? arr[5521] : arr[5520];
wire r1_2762;
assign r1_2762 = in[0]? arr[5523] : arr[5522];
wire r1_2763;
assign r1_2763 = in[0]? arr[5525] : arr[5524];
wire r1_2764;
assign r1_2764 = in[0]? arr[5527] : arr[5526];
wire r1_2765;
assign r1_2765 = in[0]? arr[5529] : arr[5528];
wire r1_2766;
assign r1_2766 = in[0]? arr[5531] : arr[5530];
wire r1_2767;
assign r1_2767 = in[0]? arr[5533] : arr[5532];
wire r1_2768;
assign r1_2768 = in[0]? arr[5535] : arr[5534];
wire r1_2769;
assign r1_2769 = in[0]? arr[5537] : arr[5536];
wire r1_2770;
assign r1_2770 = in[0]? arr[5539] : arr[5538];
wire r1_2771;
assign r1_2771 = in[0]? arr[5541] : arr[5540];
wire r1_2772;
assign r1_2772 = in[0]? arr[5543] : arr[5542];
wire r1_2773;
assign r1_2773 = in[0]? arr[5545] : arr[5544];
wire r1_2774;
assign r1_2774 = in[0]? arr[5547] : arr[5546];
wire r1_2775;
assign r1_2775 = in[0]? arr[5549] : arr[5548];
wire r1_2776;
assign r1_2776 = in[0]? arr[5551] : arr[5550];
wire r1_2777;
assign r1_2777 = in[0]? arr[5553] : arr[5552];
wire r1_2778;
assign r1_2778 = in[0]? arr[5555] : arr[5554];
wire r1_2779;
assign r1_2779 = in[0]? arr[5557] : arr[5556];
wire r1_2780;
assign r1_2780 = in[0]? arr[5559] : arr[5558];
wire r1_2781;
assign r1_2781 = in[0]? arr[5561] : arr[5560];
wire r1_2782;
assign r1_2782 = in[0]? arr[5563] : arr[5562];
wire r1_2783;
assign r1_2783 = in[0]? arr[5565] : arr[5564];
wire r1_2784;
assign r1_2784 = in[0]? arr[5567] : arr[5566];
wire r1_2785;
assign r1_2785 = in[0]? arr[5569] : arr[5568];
wire r1_2786;
assign r1_2786 = in[0]? arr[5571] : arr[5570];
wire r1_2787;
assign r1_2787 = in[0]? arr[5573] : arr[5572];
wire r1_2788;
assign r1_2788 = in[0]? arr[5575] : arr[5574];
wire r1_2789;
assign r1_2789 = in[0]? arr[5577] : arr[5576];
wire r1_2790;
assign r1_2790 = in[0]? arr[5579] : arr[5578];
wire r1_2791;
assign r1_2791 = in[0]? arr[5581] : arr[5580];
wire r1_2792;
assign r1_2792 = in[0]? arr[5583] : arr[5582];
wire r1_2793;
assign r1_2793 = in[0]? arr[5585] : arr[5584];
wire r1_2794;
assign r1_2794 = in[0]? arr[5587] : arr[5586];
wire r1_2795;
assign r1_2795 = in[0]? arr[5589] : arr[5588];
wire r1_2796;
assign r1_2796 = in[0]? arr[5591] : arr[5590];
wire r1_2797;
assign r1_2797 = in[0]? arr[5593] : arr[5592];
wire r1_2798;
assign r1_2798 = in[0]? arr[5595] : arr[5594];
wire r1_2799;
assign r1_2799 = in[0]? arr[5597] : arr[5596];
wire r1_2800;
assign r1_2800 = in[0]? arr[5599] : arr[5598];
wire r1_2801;
assign r1_2801 = in[0]? arr[5601] : arr[5600];
wire r1_2802;
assign r1_2802 = in[0]? arr[5603] : arr[5602];
wire r1_2803;
assign r1_2803 = in[0]? arr[5605] : arr[5604];
wire r1_2804;
assign r1_2804 = in[0]? arr[5607] : arr[5606];
wire r1_2805;
assign r1_2805 = in[0]? arr[5609] : arr[5608];
wire r1_2806;
assign r1_2806 = in[0]? arr[5611] : arr[5610];
wire r1_2807;
assign r1_2807 = in[0]? arr[5613] : arr[5612];
wire r1_2808;
assign r1_2808 = in[0]? arr[5615] : arr[5614];
wire r1_2809;
assign r1_2809 = in[0]? arr[5617] : arr[5616];
wire r1_2810;
assign r1_2810 = in[0]? arr[5619] : arr[5618];
wire r1_2811;
assign r1_2811 = in[0]? arr[5621] : arr[5620];
wire r1_2812;
assign r1_2812 = in[0]? arr[5623] : arr[5622];
wire r1_2813;
assign r1_2813 = in[0]? arr[5625] : arr[5624];
wire r1_2814;
assign r1_2814 = in[0]? arr[5627] : arr[5626];
wire r1_2815;
assign r1_2815 = in[0]? arr[5629] : arr[5628];
wire r1_2816;
assign r1_2816 = in[0]? arr[5631] : arr[5630];
wire r1_2817;
assign r1_2817 = in[0]? arr[5633] : arr[5632];
wire r1_2818;
assign r1_2818 = in[0]? arr[5635] : arr[5634];
wire r1_2819;
assign r1_2819 = in[0]? arr[5637] : arr[5636];
wire r1_2820;
assign r1_2820 = in[0]? arr[5639] : arr[5638];
wire r1_2821;
assign r1_2821 = in[0]? arr[5641] : arr[5640];
wire r1_2822;
assign r1_2822 = in[0]? arr[5643] : arr[5642];
wire r1_2823;
assign r1_2823 = in[0]? arr[5645] : arr[5644];
wire r1_2824;
assign r1_2824 = in[0]? arr[5647] : arr[5646];
wire r1_2825;
assign r1_2825 = in[0]? arr[5649] : arr[5648];
wire r1_2826;
assign r1_2826 = in[0]? arr[5651] : arr[5650];
wire r1_2827;
assign r1_2827 = in[0]? arr[5653] : arr[5652];
wire r1_2828;
assign r1_2828 = in[0]? arr[5655] : arr[5654];
wire r1_2829;
assign r1_2829 = in[0]? arr[5657] : arr[5656];
wire r1_2830;
assign r1_2830 = in[0]? arr[5659] : arr[5658];
wire r1_2831;
assign r1_2831 = in[0]? arr[5661] : arr[5660];
wire r1_2832;
assign r1_2832 = in[0]? arr[5663] : arr[5662];
wire r1_2833;
assign r1_2833 = in[0]? arr[5665] : arr[5664];
wire r1_2834;
assign r1_2834 = in[0]? arr[5667] : arr[5666];
wire r1_2835;
assign r1_2835 = in[0]? arr[5669] : arr[5668];
wire r1_2836;
assign r1_2836 = in[0]? arr[5671] : arr[5670];
wire r1_2837;
assign r1_2837 = in[0]? arr[5673] : arr[5672];
wire r1_2838;
assign r1_2838 = in[0]? arr[5675] : arr[5674];
wire r1_2839;
assign r1_2839 = in[0]? arr[5677] : arr[5676];
wire r1_2840;
assign r1_2840 = in[0]? arr[5679] : arr[5678];
wire r1_2841;
assign r1_2841 = in[0]? arr[5681] : arr[5680];
wire r1_2842;
assign r1_2842 = in[0]? arr[5683] : arr[5682];
wire r1_2843;
assign r1_2843 = in[0]? arr[5685] : arr[5684];
wire r1_2844;
assign r1_2844 = in[0]? arr[5687] : arr[5686];
wire r1_2845;
assign r1_2845 = in[0]? arr[5689] : arr[5688];
wire r1_2846;
assign r1_2846 = in[0]? arr[5691] : arr[5690];
wire r1_2847;
assign r1_2847 = in[0]? arr[5693] : arr[5692];
wire r1_2848;
assign r1_2848 = in[0]? arr[5695] : arr[5694];
wire r1_2849;
assign r1_2849 = in[0]? arr[5697] : arr[5696];
wire r1_2850;
assign r1_2850 = in[0]? arr[5699] : arr[5698];
wire r1_2851;
assign r1_2851 = in[0]? arr[5701] : arr[5700];
wire r1_2852;
assign r1_2852 = in[0]? arr[5703] : arr[5702];
wire r1_2853;
assign r1_2853 = in[0]? arr[5705] : arr[5704];
wire r1_2854;
assign r1_2854 = in[0]? arr[5707] : arr[5706];
wire r1_2855;
assign r1_2855 = in[0]? arr[5709] : arr[5708];
wire r1_2856;
assign r1_2856 = in[0]? arr[5711] : arr[5710];
wire r1_2857;
assign r1_2857 = in[0]? arr[5713] : arr[5712];
wire r1_2858;
assign r1_2858 = in[0]? arr[5715] : arr[5714];
wire r1_2859;
assign r1_2859 = in[0]? arr[5717] : arr[5716];
wire r1_2860;
assign r1_2860 = in[0]? arr[5719] : arr[5718];
wire r1_2861;
assign r1_2861 = in[0]? arr[5721] : arr[5720];
wire r1_2862;
assign r1_2862 = in[0]? arr[5723] : arr[5722];
wire r1_2863;
assign r1_2863 = in[0]? arr[5725] : arr[5724];
wire r1_2864;
assign r1_2864 = in[0]? arr[5727] : arr[5726];
wire r1_2865;
assign r1_2865 = in[0]? arr[5729] : arr[5728];
wire r1_2866;
assign r1_2866 = in[0]? arr[5731] : arr[5730];
wire r1_2867;
assign r1_2867 = in[0]? arr[5733] : arr[5732];
wire r1_2868;
assign r1_2868 = in[0]? arr[5735] : arr[5734];
wire r1_2869;
assign r1_2869 = in[0]? arr[5737] : arr[5736];
wire r1_2870;
assign r1_2870 = in[0]? arr[5739] : arr[5738];
wire r1_2871;
assign r1_2871 = in[0]? arr[5741] : arr[5740];
wire r1_2872;
assign r1_2872 = in[0]? arr[5743] : arr[5742];
wire r1_2873;
assign r1_2873 = in[0]? arr[5745] : arr[5744];
wire r1_2874;
assign r1_2874 = in[0]? arr[5747] : arr[5746];
wire r1_2875;
assign r1_2875 = in[0]? arr[5749] : arr[5748];
wire r1_2876;
assign r1_2876 = in[0]? arr[5751] : arr[5750];
wire r1_2877;
assign r1_2877 = in[0]? arr[5753] : arr[5752];
wire r1_2878;
assign r1_2878 = in[0]? arr[5755] : arr[5754];
wire r1_2879;
assign r1_2879 = in[0]? arr[5757] : arr[5756];
wire r1_2880;
assign r1_2880 = in[0]? arr[5759] : arr[5758];
wire r1_2881;
assign r1_2881 = in[0]? arr[5761] : arr[5760];
wire r1_2882;
assign r1_2882 = in[0]? arr[5763] : arr[5762];
wire r1_2883;
assign r1_2883 = in[0]? arr[5765] : arr[5764];
wire r1_2884;
assign r1_2884 = in[0]? arr[5767] : arr[5766];
wire r1_2885;
assign r1_2885 = in[0]? arr[5769] : arr[5768];
wire r1_2886;
assign r1_2886 = in[0]? arr[5771] : arr[5770];
wire r1_2887;
assign r1_2887 = in[0]? arr[5773] : arr[5772];
wire r1_2888;
assign r1_2888 = in[0]? arr[5775] : arr[5774];
wire r1_2889;
assign r1_2889 = in[0]? arr[5777] : arr[5776];
wire r1_2890;
assign r1_2890 = in[0]? arr[5779] : arr[5778];
wire r1_2891;
assign r1_2891 = in[0]? arr[5781] : arr[5780];
wire r1_2892;
assign r1_2892 = in[0]? arr[5783] : arr[5782];
wire r1_2893;
assign r1_2893 = in[0]? arr[5785] : arr[5784];
wire r1_2894;
assign r1_2894 = in[0]? arr[5787] : arr[5786];
wire r1_2895;
assign r1_2895 = in[0]? arr[5789] : arr[5788];
wire r1_2896;
assign r1_2896 = in[0]? arr[5791] : arr[5790];
wire r1_2897;
assign r1_2897 = in[0]? arr[5793] : arr[5792];
wire r1_2898;
assign r1_2898 = in[0]? arr[5795] : arr[5794];
wire r1_2899;
assign r1_2899 = in[0]? arr[5797] : arr[5796];
wire r1_2900;
assign r1_2900 = in[0]? arr[5799] : arr[5798];
wire r1_2901;
assign r1_2901 = in[0]? arr[5801] : arr[5800];
wire r1_2902;
assign r1_2902 = in[0]? arr[5803] : arr[5802];
wire r1_2903;
assign r1_2903 = in[0]? arr[5805] : arr[5804];
wire r1_2904;
assign r1_2904 = in[0]? arr[5807] : arr[5806];
wire r1_2905;
assign r1_2905 = in[0]? arr[5809] : arr[5808];
wire r1_2906;
assign r1_2906 = in[0]? arr[5811] : arr[5810];
wire r1_2907;
assign r1_2907 = in[0]? arr[5813] : arr[5812];
wire r1_2908;
assign r1_2908 = in[0]? arr[5815] : arr[5814];
wire r1_2909;
assign r1_2909 = in[0]? arr[5817] : arr[5816];
wire r1_2910;
assign r1_2910 = in[0]? arr[5819] : arr[5818];
wire r1_2911;
assign r1_2911 = in[0]? arr[5821] : arr[5820];
wire r1_2912;
assign r1_2912 = in[0]? arr[5823] : arr[5822];
wire r1_2913;
assign r1_2913 = in[0]? arr[5825] : arr[5824];
wire r1_2914;
assign r1_2914 = in[0]? arr[5827] : arr[5826];
wire r1_2915;
assign r1_2915 = in[0]? arr[5829] : arr[5828];
wire r1_2916;
assign r1_2916 = in[0]? arr[5831] : arr[5830];
wire r1_2917;
assign r1_2917 = in[0]? arr[5833] : arr[5832];
wire r1_2918;
assign r1_2918 = in[0]? arr[5835] : arr[5834];
wire r1_2919;
assign r1_2919 = in[0]? arr[5837] : arr[5836];
wire r1_2920;
assign r1_2920 = in[0]? arr[5839] : arr[5838];
wire r1_2921;
assign r1_2921 = in[0]? arr[5841] : arr[5840];
wire r1_2922;
assign r1_2922 = in[0]? arr[5843] : arr[5842];
wire r1_2923;
assign r1_2923 = in[0]? arr[5845] : arr[5844];
wire r1_2924;
assign r1_2924 = in[0]? arr[5847] : arr[5846];
wire r1_2925;
assign r1_2925 = in[0]? arr[5849] : arr[5848];
wire r1_2926;
assign r1_2926 = in[0]? arr[5851] : arr[5850];
wire r1_2927;
assign r1_2927 = in[0]? arr[5853] : arr[5852];
wire r1_2928;
assign r1_2928 = in[0]? arr[5855] : arr[5854];
wire r1_2929;
assign r1_2929 = in[0]? arr[5857] : arr[5856];
wire r1_2930;
assign r1_2930 = in[0]? arr[5859] : arr[5858];
wire r1_2931;
assign r1_2931 = in[0]? arr[5861] : arr[5860];
wire r1_2932;
assign r1_2932 = in[0]? arr[5863] : arr[5862];
wire r1_2933;
assign r1_2933 = in[0]? arr[5865] : arr[5864];
wire r1_2934;
assign r1_2934 = in[0]? arr[5867] : arr[5866];
wire r1_2935;
assign r1_2935 = in[0]? arr[5869] : arr[5868];
wire r1_2936;
assign r1_2936 = in[0]? arr[5871] : arr[5870];
wire r1_2937;
assign r1_2937 = in[0]? arr[5873] : arr[5872];
wire r1_2938;
assign r1_2938 = in[0]? arr[5875] : arr[5874];
wire r1_2939;
assign r1_2939 = in[0]? arr[5877] : arr[5876];
wire r1_2940;
assign r1_2940 = in[0]? arr[5879] : arr[5878];
wire r1_2941;
assign r1_2941 = in[0]? arr[5881] : arr[5880];
wire r1_2942;
assign r1_2942 = in[0]? arr[5883] : arr[5882];
wire r1_2943;
assign r1_2943 = in[0]? arr[5885] : arr[5884];
wire r1_2944;
assign r1_2944 = in[0]? arr[5887] : arr[5886];
wire r1_2945;
assign r1_2945 = in[0]? arr[5889] : arr[5888];
wire r1_2946;
assign r1_2946 = in[0]? arr[5891] : arr[5890];
wire r1_2947;
assign r1_2947 = in[0]? arr[5893] : arr[5892];
wire r1_2948;
assign r1_2948 = in[0]? arr[5895] : arr[5894];
wire r1_2949;
assign r1_2949 = in[0]? arr[5897] : arr[5896];
wire r1_2950;
assign r1_2950 = in[0]? arr[5899] : arr[5898];
wire r1_2951;
assign r1_2951 = in[0]? arr[5901] : arr[5900];
wire r1_2952;
assign r1_2952 = in[0]? arr[5903] : arr[5902];
wire r1_2953;
assign r1_2953 = in[0]? arr[5905] : arr[5904];
wire r1_2954;
assign r1_2954 = in[0]? arr[5907] : arr[5906];
wire r1_2955;
assign r1_2955 = in[0]? arr[5909] : arr[5908];
wire r1_2956;
assign r1_2956 = in[0]? arr[5911] : arr[5910];
wire r1_2957;
assign r1_2957 = in[0]? arr[5913] : arr[5912];
wire r1_2958;
assign r1_2958 = in[0]? arr[5915] : arr[5914];
wire r1_2959;
assign r1_2959 = in[0]? arr[5917] : arr[5916];
wire r1_2960;
assign r1_2960 = in[0]? arr[5919] : arr[5918];
wire r1_2961;
assign r1_2961 = in[0]? arr[5921] : arr[5920];
wire r1_2962;
assign r1_2962 = in[0]? arr[5923] : arr[5922];
wire r1_2963;
assign r1_2963 = in[0]? arr[5925] : arr[5924];
wire r1_2964;
assign r1_2964 = in[0]? arr[5927] : arr[5926];
wire r1_2965;
assign r1_2965 = in[0]? arr[5929] : arr[5928];
wire r1_2966;
assign r1_2966 = in[0]? arr[5931] : arr[5930];
wire r1_2967;
assign r1_2967 = in[0]? arr[5933] : arr[5932];
wire r1_2968;
assign r1_2968 = in[0]? arr[5935] : arr[5934];
wire r1_2969;
assign r1_2969 = in[0]? arr[5937] : arr[5936];
wire r1_2970;
assign r1_2970 = in[0]? arr[5939] : arr[5938];
wire r1_2971;
assign r1_2971 = in[0]? arr[5941] : arr[5940];
wire r1_2972;
assign r1_2972 = in[0]? arr[5943] : arr[5942];
wire r1_2973;
assign r1_2973 = in[0]? arr[5945] : arr[5944];
wire r1_2974;
assign r1_2974 = in[0]? arr[5947] : arr[5946];
wire r1_2975;
assign r1_2975 = in[0]? arr[5949] : arr[5948];
wire r1_2976;
assign r1_2976 = in[0]? arr[5951] : arr[5950];
wire r1_2977;
assign r1_2977 = in[0]? arr[5953] : arr[5952];
wire r1_2978;
assign r1_2978 = in[0]? arr[5955] : arr[5954];
wire r1_2979;
assign r1_2979 = in[0]? arr[5957] : arr[5956];
wire r1_2980;
assign r1_2980 = in[0]? arr[5959] : arr[5958];
wire r1_2981;
assign r1_2981 = in[0]? arr[5961] : arr[5960];
wire r1_2982;
assign r1_2982 = in[0]? arr[5963] : arr[5962];
wire r1_2983;
assign r1_2983 = in[0]? arr[5965] : arr[5964];
wire r1_2984;
assign r1_2984 = in[0]? arr[5967] : arr[5966];
wire r1_2985;
assign r1_2985 = in[0]? arr[5969] : arr[5968];
wire r1_2986;
assign r1_2986 = in[0]? arr[5971] : arr[5970];
wire r1_2987;
assign r1_2987 = in[0]? arr[5973] : arr[5972];
wire r1_2988;
assign r1_2988 = in[0]? arr[5975] : arr[5974];
wire r1_2989;
assign r1_2989 = in[0]? arr[5977] : arr[5976];
wire r1_2990;
assign r1_2990 = in[0]? arr[5979] : arr[5978];
wire r1_2991;
assign r1_2991 = in[0]? arr[5981] : arr[5980];
wire r1_2992;
assign r1_2992 = in[0]? arr[5983] : arr[5982];
wire r1_2993;
assign r1_2993 = in[0]? arr[5985] : arr[5984];
wire r1_2994;
assign r1_2994 = in[0]? arr[5987] : arr[5986];
wire r1_2995;
assign r1_2995 = in[0]? arr[5989] : arr[5988];
wire r1_2996;
assign r1_2996 = in[0]? arr[5991] : arr[5990];
wire r1_2997;
assign r1_2997 = in[0]? arr[5993] : arr[5992];
wire r1_2998;
assign r1_2998 = in[0]? arr[5995] : arr[5994];
wire r1_2999;
assign r1_2999 = in[0]? arr[5997] : arr[5996];
wire r1_3000;
assign r1_3000 = in[0]? arr[5999] : arr[5998];
wire r1_3001;
assign r1_3001 = in[0]? arr[6001] : arr[6000];
wire r1_3002;
assign r1_3002 = in[0]? arr[6003] : arr[6002];
wire r1_3003;
assign r1_3003 = in[0]? arr[6005] : arr[6004];
wire r1_3004;
assign r1_3004 = in[0]? arr[6007] : arr[6006];
wire r1_3005;
assign r1_3005 = in[0]? arr[6009] : arr[6008];
wire r1_3006;
assign r1_3006 = in[0]? arr[6011] : arr[6010];
wire r1_3007;
assign r1_3007 = in[0]? arr[6013] : arr[6012];
wire r1_3008;
assign r1_3008 = in[0]? arr[6015] : arr[6014];
wire r1_3009;
assign r1_3009 = in[0]? arr[6017] : arr[6016];
wire r1_3010;
assign r1_3010 = in[0]? arr[6019] : arr[6018];
wire r1_3011;
assign r1_3011 = in[0]? arr[6021] : arr[6020];
wire r1_3012;
assign r1_3012 = in[0]? arr[6023] : arr[6022];
wire r1_3013;
assign r1_3013 = in[0]? arr[6025] : arr[6024];
wire r1_3014;
assign r1_3014 = in[0]? arr[6027] : arr[6026];
wire r1_3015;
assign r1_3015 = in[0]? arr[6029] : arr[6028];
wire r1_3016;
assign r1_3016 = in[0]? arr[6031] : arr[6030];
wire r1_3017;
assign r1_3017 = in[0]? arr[6033] : arr[6032];
wire r1_3018;
assign r1_3018 = in[0]? arr[6035] : arr[6034];
wire r1_3019;
assign r1_3019 = in[0]? arr[6037] : arr[6036];
wire r1_3020;
assign r1_3020 = in[0]? arr[6039] : arr[6038];
wire r1_3021;
assign r1_3021 = in[0]? arr[6041] : arr[6040];
wire r1_3022;
assign r1_3022 = in[0]? arr[6043] : arr[6042];
wire r1_3023;
assign r1_3023 = in[0]? arr[6045] : arr[6044];
wire r1_3024;
assign r1_3024 = in[0]? arr[6047] : arr[6046];
wire r1_3025;
assign r1_3025 = in[0]? arr[6049] : arr[6048];
wire r1_3026;
assign r1_3026 = in[0]? arr[6051] : arr[6050];
wire r1_3027;
assign r1_3027 = in[0]? arr[6053] : arr[6052];
wire r1_3028;
assign r1_3028 = in[0]? arr[6055] : arr[6054];
wire r1_3029;
assign r1_3029 = in[0]? arr[6057] : arr[6056];
wire r1_3030;
assign r1_3030 = in[0]? arr[6059] : arr[6058];
wire r1_3031;
assign r1_3031 = in[0]? arr[6061] : arr[6060];
wire r1_3032;
assign r1_3032 = in[0]? arr[6063] : arr[6062];
wire r1_3033;
assign r1_3033 = in[0]? arr[6065] : arr[6064];
wire r1_3034;
assign r1_3034 = in[0]? arr[6067] : arr[6066];
wire r1_3035;
assign r1_3035 = in[0]? arr[6069] : arr[6068];
wire r1_3036;
assign r1_3036 = in[0]? arr[6071] : arr[6070];
wire r1_3037;
assign r1_3037 = in[0]? arr[6073] : arr[6072];
wire r1_3038;
assign r1_3038 = in[0]? arr[6075] : arr[6074];
wire r1_3039;
assign r1_3039 = in[0]? arr[6077] : arr[6076];
wire r1_3040;
assign r1_3040 = in[0]? arr[6079] : arr[6078];
wire r1_3041;
assign r1_3041 = in[0]? arr[6081] : arr[6080];
wire r1_3042;
assign r1_3042 = in[0]? arr[6083] : arr[6082];
wire r1_3043;
assign r1_3043 = in[0]? arr[6085] : arr[6084];
wire r1_3044;
assign r1_3044 = in[0]? arr[6087] : arr[6086];
wire r1_3045;
assign r1_3045 = in[0]? arr[6089] : arr[6088];
wire r1_3046;
assign r1_3046 = in[0]? arr[6091] : arr[6090];
wire r1_3047;
assign r1_3047 = in[0]? arr[6093] : arr[6092];
wire r1_3048;
assign r1_3048 = in[0]? arr[6095] : arr[6094];
wire r1_3049;
assign r1_3049 = in[0]? arr[6097] : arr[6096];
wire r1_3050;
assign r1_3050 = in[0]? arr[6099] : arr[6098];
wire r1_3051;
assign r1_3051 = in[0]? arr[6101] : arr[6100];
wire r1_3052;
assign r1_3052 = in[0]? arr[6103] : arr[6102];
wire r1_3053;
assign r1_3053 = in[0]? arr[6105] : arr[6104];
wire r1_3054;
assign r1_3054 = in[0]? arr[6107] : arr[6106];
wire r1_3055;
assign r1_3055 = in[0]? arr[6109] : arr[6108];
wire r1_3056;
assign r1_3056 = in[0]? arr[6111] : arr[6110];
wire r1_3057;
assign r1_3057 = in[0]? arr[6113] : arr[6112];
wire r1_3058;
assign r1_3058 = in[0]? arr[6115] : arr[6114];
wire r1_3059;
assign r1_3059 = in[0]? arr[6117] : arr[6116];
wire r1_3060;
assign r1_3060 = in[0]? arr[6119] : arr[6118];
wire r1_3061;
assign r1_3061 = in[0]? arr[6121] : arr[6120];
wire r1_3062;
assign r1_3062 = in[0]? arr[6123] : arr[6122];
wire r1_3063;
assign r1_3063 = in[0]? arr[6125] : arr[6124];
wire r1_3064;
assign r1_3064 = in[0]? arr[6127] : arr[6126];
wire r1_3065;
assign r1_3065 = in[0]? arr[6129] : arr[6128];
wire r1_3066;
assign r1_3066 = in[0]? arr[6131] : arr[6130];
wire r1_3067;
assign r1_3067 = in[0]? arr[6133] : arr[6132];
wire r1_3068;
assign r1_3068 = in[0]? arr[6135] : arr[6134];
wire r1_3069;
assign r1_3069 = in[0]? arr[6137] : arr[6136];
wire r1_3070;
assign r1_3070 = in[0]? arr[6139] : arr[6138];
wire r1_3071;
assign r1_3071 = in[0]? arr[6141] : arr[6140];
wire r1_3072;
assign r1_3072 = in[0]? arr[6143] : arr[6142];
wire r2_1;
assign r2_1 = in[1]? r1_2 : r1_1;
wire r2_2;
assign r2_2 = in[1]? r1_4 : r1_3;
wire r2_3;
assign r2_3 = in[1]? r1_6 : r1_5;
wire r2_4;
assign r2_4 = in[1]? r1_8 : r1_7;
wire r2_5;
assign r2_5 = in[1]? r1_10 : r1_9;
wire r2_6;
assign r2_6 = in[1]? r1_12 : r1_11;
wire r2_7;
assign r2_7 = in[1]? r1_14 : r1_13;
wire r2_8;
assign r2_8 = in[1]? r1_16 : r1_15;
wire r2_9;
assign r2_9 = in[1]? r1_18 : r1_17;
wire r2_10;
assign r2_10 = in[1]? r1_20 : r1_19;
wire r2_11;
assign r2_11 = in[1]? r1_22 : r1_21;
wire r2_12;
assign r2_12 = in[1]? r1_24 : r1_23;
wire r2_13;
assign r2_13 = in[1]? r1_26 : r1_25;
wire r2_14;
assign r2_14 = in[1]? r1_28 : r1_27;
wire r2_15;
assign r2_15 = in[1]? r1_30 : r1_29;
wire r2_16;
assign r2_16 = in[1]? r1_32 : r1_31;
wire r2_17;
assign r2_17 = in[1]? r1_34 : r1_33;
wire r2_18;
assign r2_18 = in[1]? r1_36 : r1_35;
wire r2_19;
assign r2_19 = in[1]? r1_38 : r1_37;
wire r2_20;
assign r2_20 = in[1]? r1_40 : r1_39;
wire r2_21;
assign r2_21 = in[1]? r1_42 : r1_41;
wire r2_22;
assign r2_22 = in[1]? r1_44 : r1_43;
wire r2_23;
assign r2_23 = in[1]? r1_46 : r1_45;
wire r2_24;
assign r2_24 = in[1]? r1_48 : r1_47;
wire r2_25;
assign r2_25 = in[1]? r1_50 : r1_49;
wire r2_26;
assign r2_26 = in[1]? r1_52 : r1_51;
wire r2_27;
assign r2_27 = in[1]? r1_54 : r1_53;
wire r2_28;
assign r2_28 = in[1]? r1_56 : r1_55;
wire r2_29;
assign r2_29 = in[1]? r1_58 : r1_57;
wire r2_30;
assign r2_30 = in[1]? r1_60 : r1_59;
wire r2_31;
assign r2_31 = in[1]? r1_62 : r1_61;
wire r2_32;
assign r2_32 = in[1]? r1_64 : r1_63;
wire r2_33;
assign r2_33 = in[1]? r1_66 : r1_65;
wire r2_34;
assign r2_34 = in[1]? r1_68 : r1_67;
wire r2_35;
assign r2_35 = in[1]? r1_70 : r1_69;
wire r2_36;
assign r2_36 = in[1]? r1_72 : r1_71;
wire r2_37;
assign r2_37 = in[1]? r1_74 : r1_73;
wire r2_38;
assign r2_38 = in[1]? r1_76 : r1_75;
wire r2_39;
assign r2_39 = in[1]? r1_78 : r1_77;
wire r2_40;
assign r2_40 = in[1]? r1_80 : r1_79;
wire r2_41;
assign r2_41 = in[1]? r1_82 : r1_81;
wire r2_42;
assign r2_42 = in[1]? r1_84 : r1_83;
wire r2_43;
assign r2_43 = in[1]? r1_86 : r1_85;
wire r2_44;
assign r2_44 = in[1]? r1_88 : r1_87;
wire r2_45;
assign r2_45 = in[1]? r1_90 : r1_89;
wire r2_46;
assign r2_46 = in[1]? r1_92 : r1_91;
wire r2_47;
assign r2_47 = in[1]? r1_94 : r1_93;
wire r2_48;
assign r2_48 = in[1]? r1_96 : r1_95;
wire r2_49;
assign r2_49 = in[1]? r1_98 : r1_97;
wire r2_50;
assign r2_50 = in[1]? r1_100 : r1_99;
wire r2_51;
assign r2_51 = in[1]? r1_102 : r1_101;
wire r2_52;
assign r2_52 = in[1]? r1_104 : r1_103;
wire r2_53;
assign r2_53 = in[1]? r1_106 : r1_105;
wire r2_54;
assign r2_54 = in[1]? r1_108 : r1_107;
wire r2_55;
assign r2_55 = in[1]? r1_110 : r1_109;
wire r2_56;
assign r2_56 = in[1]? r1_112 : r1_111;
wire r2_57;
assign r2_57 = in[1]? r1_114 : r1_113;
wire r2_58;
assign r2_58 = in[1]? r1_116 : r1_115;
wire r2_59;
assign r2_59 = in[1]? r1_118 : r1_117;
wire r2_60;
assign r2_60 = in[1]? r1_120 : r1_119;
wire r2_61;
assign r2_61 = in[1]? r1_122 : r1_121;
wire r2_62;
assign r2_62 = in[1]? r1_124 : r1_123;
wire r2_63;
assign r2_63 = in[1]? r1_126 : r1_125;
wire r2_64;
assign r2_64 = in[1]? r1_128 : r1_127;
wire r2_65;
assign r2_65 = in[1]? r1_130 : r1_129;
wire r2_66;
assign r2_66 = in[1]? r1_132 : r1_131;
wire r2_67;
assign r2_67 = in[1]? r1_134 : r1_133;
wire r2_68;
assign r2_68 = in[1]? r1_136 : r1_135;
wire r2_69;
assign r2_69 = in[1]? r1_138 : r1_137;
wire r2_70;
assign r2_70 = in[1]? r1_140 : r1_139;
wire r2_71;
assign r2_71 = in[1]? r1_142 : r1_141;
wire r2_72;
assign r2_72 = in[1]? r1_144 : r1_143;
wire r2_73;
assign r2_73 = in[1]? r1_146 : r1_145;
wire r2_74;
assign r2_74 = in[1]? r1_148 : r1_147;
wire r2_75;
assign r2_75 = in[1]? r1_150 : r1_149;
wire r2_76;
assign r2_76 = in[1]? r1_152 : r1_151;
wire r2_77;
assign r2_77 = in[1]? r1_154 : r1_153;
wire r2_78;
assign r2_78 = in[1]? r1_156 : r1_155;
wire r2_79;
assign r2_79 = in[1]? r1_158 : r1_157;
wire r2_80;
assign r2_80 = in[1]? r1_160 : r1_159;
wire r2_81;
assign r2_81 = in[1]? r1_162 : r1_161;
wire r2_82;
assign r2_82 = in[1]? r1_164 : r1_163;
wire r2_83;
assign r2_83 = in[1]? r1_166 : r1_165;
wire r2_84;
assign r2_84 = in[1]? r1_168 : r1_167;
wire r2_85;
assign r2_85 = in[1]? r1_170 : r1_169;
wire r2_86;
assign r2_86 = in[1]? r1_172 : r1_171;
wire r2_87;
assign r2_87 = in[1]? r1_174 : r1_173;
wire r2_88;
assign r2_88 = in[1]? r1_176 : r1_175;
wire r2_89;
assign r2_89 = in[1]? r1_178 : r1_177;
wire r2_90;
assign r2_90 = in[1]? r1_180 : r1_179;
wire r2_91;
assign r2_91 = in[1]? r1_182 : r1_181;
wire r2_92;
assign r2_92 = in[1]? r1_184 : r1_183;
wire r2_93;
assign r2_93 = in[1]? r1_186 : r1_185;
wire r2_94;
assign r2_94 = in[1]? r1_188 : r1_187;
wire r2_95;
assign r2_95 = in[1]? r1_190 : r1_189;
wire r2_96;
assign r2_96 = in[1]? r1_192 : r1_191;
wire r2_97;
assign r2_97 = in[1]? r1_194 : r1_193;
wire r2_98;
assign r2_98 = in[1]? r1_196 : r1_195;
wire r2_99;
assign r2_99 = in[1]? r1_198 : r1_197;
wire r2_100;
assign r2_100 = in[1]? r1_200 : r1_199;
wire r2_101;
assign r2_101 = in[1]? r1_202 : r1_201;
wire r2_102;
assign r2_102 = in[1]? r1_204 : r1_203;
wire r2_103;
assign r2_103 = in[1]? r1_206 : r1_205;
wire r2_104;
assign r2_104 = in[1]? r1_208 : r1_207;
wire r2_105;
assign r2_105 = in[1]? r1_210 : r1_209;
wire r2_106;
assign r2_106 = in[1]? r1_212 : r1_211;
wire r2_107;
assign r2_107 = in[1]? r1_214 : r1_213;
wire r2_108;
assign r2_108 = in[1]? r1_216 : r1_215;
wire r2_109;
assign r2_109 = in[1]? r1_218 : r1_217;
wire r2_110;
assign r2_110 = in[1]? r1_220 : r1_219;
wire r2_111;
assign r2_111 = in[1]? r1_222 : r1_221;
wire r2_112;
assign r2_112 = in[1]? r1_224 : r1_223;
wire r2_113;
assign r2_113 = in[1]? r1_226 : r1_225;
wire r2_114;
assign r2_114 = in[1]? r1_228 : r1_227;
wire r2_115;
assign r2_115 = in[1]? r1_230 : r1_229;
wire r2_116;
assign r2_116 = in[1]? r1_232 : r1_231;
wire r2_117;
assign r2_117 = in[1]? r1_234 : r1_233;
wire r2_118;
assign r2_118 = in[1]? r1_236 : r1_235;
wire r2_119;
assign r2_119 = in[1]? r1_238 : r1_237;
wire r2_120;
assign r2_120 = in[1]? r1_240 : r1_239;
wire r2_121;
assign r2_121 = in[1]? r1_242 : r1_241;
wire r2_122;
assign r2_122 = in[1]? r1_244 : r1_243;
wire r2_123;
assign r2_123 = in[1]? r1_246 : r1_245;
wire r2_124;
assign r2_124 = in[1]? r1_248 : r1_247;
wire r2_125;
assign r2_125 = in[1]? r1_250 : r1_249;
wire r2_126;
assign r2_126 = in[1]? r1_252 : r1_251;
wire r2_127;
assign r2_127 = in[1]? r1_254 : r1_253;
wire r2_128;
assign r2_128 = in[1]? r1_256 : r1_255;
wire r2_129;
assign r2_129 = in[1]? r1_258 : r1_257;
wire r2_130;
assign r2_130 = in[1]? r1_260 : r1_259;
wire r2_131;
assign r2_131 = in[1]? r1_262 : r1_261;
wire r2_132;
assign r2_132 = in[1]? r1_264 : r1_263;
wire r2_133;
assign r2_133 = in[1]? r1_266 : r1_265;
wire r2_134;
assign r2_134 = in[1]? r1_268 : r1_267;
wire r2_135;
assign r2_135 = in[1]? r1_270 : r1_269;
wire r2_136;
assign r2_136 = in[1]? r1_272 : r1_271;
wire r2_137;
assign r2_137 = in[1]? r1_274 : r1_273;
wire r2_138;
assign r2_138 = in[1]? r1_276 : r1_275;
wire r2_139;
assign r2_139 = in[1]? r1_278 : r1_277;
wire r2_140;
assign r2_140 = in[1]? r1_280 : r1_279;
wire r2_141;
assign r2_141 = in[1]? r1_282 : r1_281;
wire r2_142;
assign r2_142 = in[1]? r1_284 : r1_283;
wire r2_143;
assign r2_143 = in[1]? r1_286 : r1_285;
wire r2_144;
assign r2_144 = in[1]? r1_288 : r1_287;
wire r2_145;
assign r2_145 = in[1]? r1_290 : r1_289;
wire r2_146;
assign r2_146 = in[1]? r1_292 : r1_291;
wire r2_147;
assign r2_147 = in[1]? r1_294 : r1_293;
wire r2_148;
assign r2_148 = in[1]? r1_296 : r1_295;
wire r2_149;
assign r2_149 = in[1]? r1_298 : r1_297;
wire r2_150;
assign r2_150 = in[1]? r1_300 : r1_299;
wire r2_151;
assign r2_151 = in[1]? r1_302 : r1_301;
wire r2_152;
assign r2_152 = in[1]? r1_304 : r1_303;
wire r2_153;
assign r2_153 = in[1]? r1_306 : r1_305;
wire r2_154;
assign r2_154 = in[1]? r1_308 : r1_307;
wire r2_155;
assign r2_155 = in[1]? r1_310 : r1_309;
wire r2_156;
assign r2_156 = in[1]? r1_312 : r1_311;
wire r2_157;
assign r2_157 = in[1]? r1_314 : r1_313;
wire r2_158;
assign r2_158 = in[1]? r1_316 : r1_315;
wire r2_159;
assign r2_159 = in[1]? r1_318 : r1_317;
wire r2_160;
assign r2_160 = in[1]? r1_320 : r1_319;
wire r2_161;
assign r2_161 = in[1]? r1_322 : r1_321;
wire r2_162;
assign r2_162 = in[1]? r1_324 : r1_323;
wire r2_163;
assign r2_163 = in[1]? r1_326 : r1_325;
wire r2_164;
assign r2_164 = in[1]? r1_328 : r1_327;
wire r2_165;
assign r2_165 = in[1]? r1_330 : r1_329;
wire r2_166;
assign r2_166 = in[1]? r1_332 : r1_331;
wire r2_167;
assign r2_167 = in[1]? r1_334 : r1_333;
wire r2_168;
assign r2_168 = in[1]? r1_336 : r1_335;
wire r2_169;
assign r2_169 = in[1]? r1_338 : r1_337;
wire r2_170;
assign r2_170 = in[1]? r1_340 : r1_339;
wire r2_171;
assign r2_171 = in[1]? r1_342 : r1_341;
wire r2_172;
assign r2_172 = in[1]? r1_344 : r1_343;
wire r2_173;
assign r2_173 = in[1]? r1_346 : r1_345;
wire r2_174;
assign r2_174 = in[1]? r1_348 : r1_347;
wire r2_175;
assign r2_175 = in[1]? r1_350 : r1_349;
wire r2_176;
assign r2_176 = in[1]? r1_352 : r1_351;
wire r2_177;
assign r2_177 = in[1]? r1_354 : r1_353;
wire r2_178;
assign r2_178 = in[1]? r1_356 : r1_355;
wire r2_179;
assign r2_179 = in[1]? r1_358 : r1_357;
wire r2_180;
assign r2_180 = in[1]? r1_360 : r1_359;
wire r2_181;
assign r2_181 = in[1]? r1_362 : r1_361;
wire r2_182;
assign r2_182 = in[1]? r1_364 : r1_363;
wire r2_183;
assign r2_183 = in[1]? r1_366 : r1_365;
wire r2_184;
assign r2_184 = in[1]? r1_368 : r1_367;
wire r2_185;
assign r2_185 = in[1]? r1_370 : r1_369;
wire r2_186;
assign r2_186 = in[1]? r1_372 : r1_371;
wire r2_187;
assign r2_187 = in[1]? r1_374 : r1_373;
wire r2_188;
assign r2_188 = in[1]? r1_376 : r1_375;
wire r2_189;
assign r2_189 = in[1]? r1_378 : r1_377;
wire r2_190;
assign r2_190 = in[1]? r1_380 : r1_379;
wire r2_191;
assign r2_191 = in[1]? r1_382 : r1_381;
wire r2_192;
assign r2_192 = in[1]? r1_384 : r1_383;
wire r2_193;
assign r2_193 = in[1]? r1_386 : r1_385;
wire r2_194;
assign r2_194 = in[1]? r1_388 : r1_387;
wire r2_195;
assign r2_195 = in[1]? r1_390 : r1_389;
wire r2_196;
assign r2_196 = in[1]? r1_392 : r1_391;
wire r2_197;
assign r2_197 = in[1]? r1_394 : r1_393;
wire r2_198;
assign r2_198 = in[1]? r1_396 : r1_395;
wire r2_199;
assign r2_199 = in[1]? r1_398 : r1_397;
wire r2_200;
assign r2_200 = in[1]? r1_400 : r1_399;
wire r2_201;
assign r2_201 = in[1]? r1_402 : r1_401;
wire r2_202;
assign r2_202 = in[1]? r1_404 : r1_403;
wire r2_203;
assign r2_203 = in[1]? r1_406 : r1_405;
wire r2_204;
assign r2_204 = in[1]? r1_408 : r1_407;
wire r2_205;
assign r2_205 = in[1]? r1_410 : r1_409;
wire r2_206;
assign r2_206 = in[1]? r1_412 : r1_411;
wire r2_207;
assign r2_207 = in[1]? r1_414 : r1_413;
wire r2_208;
assign r2_208 = in[1]? r1_416 : r1_415;
wire r2_209;
assign r2_209 = in[1]? r1_418 : r1_417;
wire r2_210;
assign r2_210 = in[1]? r1_420 : r1_419;
wire r2_211;
assign r2_211 = in[1]? r1_422 : r1_421;
wire r2_212;
assign r2_212 = in[1]? r1_424 : r1_423;
wire r2_213;
assign r2_213 = in[1]? r1_426 : r1_425;
wire r2_214;
assign r2_214 = in[1]? r1_428 : r1_427;
wire r2_215;
assign r2_215 = in[1]? r1_430 : r1_429;
wire r2_216;
assign r2_216 = in[1]? r1_432 : r1_431;
wire r2_217;
assign r2_217 = in[1]? r1_434 : r1_433;
wire r2_218;
assign r2_218 = in[1]? r1_436 : r1_435;
wire r2_219;
assign r2_219 = in[1]? r1_438 : r1_437;
wire r2_220;
assign r2_220 = in[1]? r1_440 : r1_439;
wire r2_221;
assign r2_221 = in[1]? r1_442 : r1_441;
wire r2_222;
assign r2_222 = in[1]? r1_444 : r1_443;
wire r2_223;
assign r2_223 = in[1]? r1_446 : r1_445;
wire r2_224;
assign r2_224 = in[1]? r1_448 : r1_447;
wire r2_225;
assign r2_225 = in[1]? r1_450 : r1_449;
wire r2_226;
assign r2_226 = in[1]? r1_452 : r1_451;
wire r2_227;
assign r2_227 = in[1]? r1_454 : r1_453;
wire r2_228;
assign r2_228 = in[1]? r1_456 : r1_455;
wire r2_229;
assign r2_229 = in[1]? r1_458 : r1_457;
wire r2_230;
assign r2_230 = in[1]? r1_460 : r1_459;
wire r2_231;
assign r2_231 = in[1]? r1_462 : r1_461;
wire r2_232;
assign r2_232 = in[1]? r1_464 : r1_463;
wire r2_233;
assign r2_233 = in[1]? r1_466 : r1_465;
wire r2_234;
assign r2_234 = in[1]? r1_468 : r1_467;
wire r2_235;
assign r2_235 = in[1]? r1_470 : r1_469;
wire r2_236;
assign r2_236 = in[1]? r1_472 : r1_471;
wire r2_237;
assign r2_237 = in[1]? r1_474 : r1_473;
wire r2_238;
assign r2_238 = in[1]? r1_476 : r1_475;
wire r2_239;
assign r2_239 = in[1]? r1_478 : r1_477;
wire r2_240;
assign r2_240 = in[1]? r1_480 : r1_479;
wire r2_241;
assign r2_241 = in[1]? r1_482 : r1_481;
wire r2_242;
assign r2_242 = in[1]? r1_484 : r1_483;
wire r2_243;
assign r2_243 = in[1]? r1_486 : r1_485;
wire r2_244;
assign r2_244 = in[1]? r1_488 : r1_487;
wire r2_245;
assign r2_245 = in[1]? r1_490 : r1_489;
wire r2_246;
assign r2_246 = in[1]? r1_492 : r1_491;
wire r2_247;
assign r2_247 = in[1]? r1_494 : r1_493;
wire r2_248;
assign r2_248 = in[1]? r1_496 : r1_495;
wire r2_249;
assign r2_249 = in[1]? r1_498 : r1_497;
wire r2_250;
assign r2_250 = in[1]? r1_500 : r1_499;
wire r2_251;
assign r2_251 = in[1]? r1_502 : r1_501;
wire r2_252;
assign r2_252 = in[1]? r1_504 : r1_503;
wire r2_253;
assign r2_253 = in[1]? r1_506 : r1_505;
wire r2_254;
assign r2_254 = in[1]? r1_508 : r1_507;
wire r2_255;
assign r2_255 = in[1]? r1_510 : r1_509;
wire r2_256;
assign r2_256 = in[1]? r1_512 : r1_511;
wire r2_257;
assign r2_257 = in[1]? r1_514 : r1_513;
wire r2_258;
assign r2_258 = in[1]? r1_516 : r1_515;
wire r2_259;
assign r2_259 = in[1]? r1_518 : r1_517;
wire r2_260;
assign r2_260 = in[1]? r1_520 : r1_519;
wire r2_261;
assign r2_261 = in[1]? r1_522 : r1_521;
wire r2_262;
assign r2_262 = in[1]? r1_524 : r1_523;
wire r2_263;
assign r2_263 = in[1]? r1_526 : r1_525;
wire r2_264;
assign r2_264 = in[1]? r1_528 : r1_527;
wire r2_265;
assign r2_265 = in[1]? r1_530 : r1_529;
wire r2_266;
assign r2_266 = in[1]? r1_532 : r1_531;
wire r2_267;
assign r2_267 = in[1]? r1_534 : r1_533;
wire r2_268;
assign r2_268 = in[1]? r1_536 : r1_535;
wire r2_269;
assign r2_269 = in[1]? r1_538 : r1_537;
wire r2_270;
assign r2_270 = in[1]? r1_540 : r1_539;
wire r2_271;
assign r2_271 = in[1]? r1_542 : r1_541;
wire r2_272;
assign r2_272 = in[1]? r1_544 : r1_543;
wire r2_273;
assign r2_273 = in[1]? r1_546 : r1_545;
wire r2_274;
assign r2_274 = in[1]? r1_548 : r1_547;
wire r2_275;
assign r2_275 = in[1]? r1_550 : r1_549;
wire r2_276;
assign r2_276 = in[1]? r1_552 : r1_551;
wire r2_277;
assign r2_277 = in[1]? r1_554 : r1_553;
wire r2_278;
assign r2_278 = in[1]? r1_556 : r1_555;
wire r2_279;
assign r2_279 = in[1]? r1_558 : r1_557;
wire r2_280;
assign r2_280 = in[1]? r1_560 : r1_559;
wire r2_281;
assign r2_281 = in[1]? r1_562 : r1_561;
wire r2_282;
assign r2_282 = in[1]? r1_564 : r1_563;
wire r2_283;
assign r2_283 = in[1]? r1_566 : r1_565;
wire r2_284;
assign r2_284 = in[1]? r1_568 : r1_567;
wire r2_285;
assign r2_285 = in[1]? r1_570 : r1_569;
wire r2_286;
assign r2_286 = in[1]? r1_572 : r1_571;
wire r2_287;
assign r2_287 = in[1]? r1_574 : r1_573;
wire r2_288;
assign r2_288 = in[1]? r1_576 : r1_575;
wire r2_289;
assign r2_289 = in[1]? r1_578 : r1_577;
wire r2_290;
assign r2_290 = in[1]? r1_580 : r1_579;
wire r2_291;
assign r2_291 = in[1]? r1_582 : r1_581;
wire r2_292;
assign r2_292 = in[1]? r1_584 : r1_583;
wire r2_293;
assign r2_293 = in[1]? r1_586 : r1_585;
wire r2_294;
assign r2_294 = in[1]? r1_588 : r1_587;
wire r2_295;
assign r2_295 = in[1]? r1_590 : r1_589;
wire r2_296;
assign r2_296 = in[1]? r1_592 : r1_591;
wire r2_297;
assign r2_297 = in[1]? r1_594 : r1_593;
wire r2_298;
assign r2_298 = in[1]? r1_596 : r1_595;
wire r2_299;
assign r2_299 = in[1]? r1_598 : r1_597;
wire r2_300;
assign r2_300 = in[1]? r1_600 : r1_599;
wire r2_301;
assign r2_301 = in[1]? r1_602 : r1_601;
wire r2_302;
assign r2_302 = in[1]? r1_604 : r1_603;
wire r2_303;
assign r2_303 = in[1]? r1_606 : r1_605;
wire r2_304;
assign r2_304 = in[1]? r1_608 : r1_607;
wire r2_305;
assign r2_305 = in[1]? r1_610 : r1_609;
wire r2_306;
assign r2_306 = in[1]? r1_612 : r1_611;
wire r2_307;
assign r2_307 = in[1]? r1_614 : r1_613;
wire r2_308;
assign r2_308 = in[1]? r1_616 : r1_615;
wire r2_309;
assign r2_309 = in[1]? r1_618 : r1_617;
wire r2_310;
assign r2_310 = in[1]? r1_620 : r1_619;
wire r2_311;
assign r2_311 = in[1]? r1_622 : r1_621;
wire r2_312;
assign r2_312 = in[1]? r1_624 : r1_623;
wire r2_313;
assign r2_313 = in[1]? r1_626 : r1_625;
wire r2_314;
assign r2_314 = in[1]? r1_628 : r1_627;
wire r2_315;
assign r2_315 = in[1]? r1_630 : r1_629;
wire r2_316;
assign r2_316 = in[1]? r1_632 : r1_631;
wire r2_317;
assign r2_317 = in[1]? r1_634 : r1_633;
wire r2_318;
assign r2_318 = in[1]? r1_636 : r1_635;
wire r2_319;
assign r2_319 = in[1]? r1_638 : r1_637;
wire r2_320;
assign r2_320 = in[1]? r1_640 : r1_639;
wire r2_321;
assign r2_321 = in[1]? r1_642 : r1_641;
wire r2_322;
assign r2_322 = in[1]? r1_644 : r1_643;
wire r2_323;
assign r2_323 = in[1]? r1_646 : r1_645;
wire r2_324;
assign r2_324 = in[1]? r1_648 : r1_647;
wire r2_325;
assign r2_325 = in[1]? r1_650 : r1_649;
wire r2_326;
assign r2_326 = in[1]? r1_652 : r1_651;
wire r2_327;
assign r2_327 = in[1]? r1_654 : r1_653;
wire r2_328;
assign r2_328 = in[1]? r1_656 : r1_655;
wire r2_329;
assign r2_329 = in[1]? r1_658 : r1_657;
wire r2_330;
assign r2_330 = in[1]? r1_660 : r1_659;
wire r2_331;
assign r2_331 = in[1]? r1_662 : r1_661;
wire r2_332;
assign r2_332 = in[1]? r1_664 : r1_663;
wire r2_333;
assign r2_333 = in[1]? r1_666 : r1_665;
wire r2_334;
assign r2_334 = in[1]? r1_668 : r1_667;
wire r2_335;
assign r2_335 = in[1]? r1_670 : r1_669;
wire r2_336;
assign r2_336 = in[1]? r1_672 : r1_671;
wire r2_337;
assign r2_337 = in[1]? r1_674 : r1_673;
wire r2_338;
assign r2_338 = in[1]? r1_676 : r1_675;
wire r2_339;
assign r2_339 = in[1]? r1_678 : r1_677;
wire r2_340;
assign r2_340 = in[1]? r1_680 : r1_679;
wire r2_341;
assign r2_341 = in[1]? r1_682 : r1_681;
wire r2_342;
assign r2_342 = in[1]? r1_684 : r1_683;
wire r2_343;
assign r2_343 = in[1]? r1_686 : r1_685;
wire r2_344;
assign r2_344 = in[1]? r1_688 : r1_687;
wire r2_345;
assign r2_345 = in[1]? r1_690 : r1_689;
wire r2_346;
assign r2_346 = in[1]? r1_692 : r1_691;
wire r2_347;
assign r2_347 = in[1]? r1_694 : r1_693;
wire r2_348;
assign r2_348 = in[1]? r1_696 : r1_695;
wire r2_349;
assign r2_349 = in[1]? r1_698 : r1_697;
wire r2_350;
assign r2_350 = in[1]? r1_700 : r1_699;
wire r2_351;
assign r2_351 = in[1]? r1_702 : r1_701;
wire r2_352;
assign r2_352 = in[1]? r1_704 : r1_703;
wire r2_353;
assign r2_353 = in[1]? r1_706 : r1_705;
wire r2_354;
assign r2_354 = in[1]? r1_708 : r1_707;
wire r2_355;
assign r2_355 = in[1]? r1_710 : r1_709;
wire r2_356;
assign r2_356 = in[1]? r1_712 : r1_711;
wire r2_357;
assign r2_357 = in[1]? r1_714 : r1_713;
wire r2_358;
assign r2_358 = in[1]? r1_716 : r1_715;
wire r2_359;
assign r2_359 = in[1]? r1_718 : r1_717;
wire r2_360;
assign r2_360 = in[1]? r1_720 : r1_719;
wire r2_361;
assign r2_361 = in[1]? r1_722 : r1_721;
wire r2_362;
assign r2_362 = in[1]? r1_724 : r1_723;
wire r2_363;
assign r2_363 = in[1]? r1_726 : r1_725;
wire r2_364;
assign r2_364 = in[1]? r1_728 : r1_727;
wire r2_365;
assign r2_365 = in[1]? r1_730 : r1_729;
wire r2_366;
assign r2_366 = in[1]? r1_732 : r1_731;
wire r2_367;
assign r2_367 = in[1]? r1_734 : r1_733;
wire r2_368;
assign r2_368 = in[1]? r1_736 : r1_735;
wire r2_369;
assign r2_369 = in[1]? r1_738 : r1_737;
wire r2_370;
assign r2_370 = in[1]? r1_740 : r1_739;
wire r2_371;
assign r2_371 = in[1]? r1_742 : r1_741;
wire r2_372;
assign r2_372 = in[1]? r1_744 : r1_743;
wire r2_373;
assign r2_373 = in[1]? r1_746 : r1_745;
wire r2_374;
assign r2_374 = in[1]? r1_748 : r1_747;
wire r2_375;
assign r2_375 = in[1]? r1_750 : r1_749;
wire r2_376;
assign r2_376 = in[1]? r1_752 : r1_751;
wire r2_377;
assign r2_377 = in[1]? r1_754 : r1_753;
wire r2_378;
assign r2_378 = in[1]? r1_756 : r1_755;
wire r2_379;
assign r2_379 = in[1]? r1_758 : r1_757;
wire r2_380;
assign r2_380 = in[1]? r1_760 : r1_759;
wire r2_381;
assign r2_381 = in[1]? r1_762 : r1_761;
wire r2_382;
assign r2_382 = in[1]? r1_764 : r1_763;
wire r2_383;
assign r2_383 = in[1]? r1_766 : r1_765;
wire r2_384;
assign r2_384 = in[1]? r1_768 : r1_767;
wire r2_385;
assign r2_385 = in[1]? r1_770 : r1_769;
wire r2_386;
assign r2_386 = in[1]? r1_772 : r1_771;
wire r2_387;
assign r2_387 = in[1]? r1_774 : r1_773;
wire r2_388;
assign r2_388 = in[1]? r1_776 : r1_775;
wire r2_389;
assign r2_389 = in[1]? r1_778 : r1_777;
wire r2_390;
assign r2_390 = in[1]? r1_780 : r1_779;
wire r2_391;
assign r2_391 = in[1]? r1_782 : r1_781;
wire r2_392;
assign r2_392 = in[1]? r1_784 : r1_783;
wire r2_393;
assign r2_393 = in[1]? r1_786 : r1_785;
wire r2_394;
assign r2_394 = in[1]? r1_788 : r1_787;
wire r2_395;
assign r2_395 = in[1]? r1_790 : r1_789;
wire r2_396;
assign r2_396 = in[1]? r1_792 : r1_791;
wire r2_397;
assign r2_397 = in[1]? r1_794 : r1_793;
wire r2_398;
assign r2_398 = in[1]? r1_796 : r1_795;
wire r2_399;
assign r2_399 = in[1]? r1_798 : r1_797;
wire r2_400;
assign r2_400 = in[1]? r1_800 : r1_799;
wire r2_401;
assign r2_401 = in[1]? r1_802 : r1_801;
wire r2_402;
assign r2_402 = in[1]? r1_804 : r1_803;
wire r2_403;
assign r2_403 = in[1]? r1_806 : r1_805;
wire r2_404;
assign r2_404 = in[1]? r1_808 : r1_807;
wire r2_405;
assign r2_405 = in[1]? r1_810 : r1_809;
wire r2_406;
assign r2_406 = in[1]? r1_812 : r1_811;
wire r2_407;
assign r2_407 = in[1]? r1_814 : r1_813;
wire r2_408;
assign r2_408 = in[1]? r1_816 : r1_815;
wire r2_409;
assign r2_409 = in[1]? r1_818 : r1_817;
wire r2_410;
assign r2_410 = in[1]? r1_820 : r1_819;
wire r2_411;
assign r2_411 = in[1]? r1_822 : r1_821;
wire r2_412;
assign r2_412 = in[1]? r1_824 : r1_823;
wire r2_413;
assign r2_413 = in[1]? r1_826 : r1_825;
wire r2_414;
assign r2_414 = in[1]? r1_828 : r1_827;
wire r2_415;
assign r2_415 = in[1]? r1_830 : r1_829;
wire r2_416;
assign r2_416 = in[1]? r1_832 : r1_831;
wire r2_417;
assign r2_417 = in[1]? r1_834 : r1_833;
wire r2_418;
assign r2_418 = in[1]? r1_836 : r1_835;
wire r2_419;
assign r2_419 = in[1]? r1_838 : r1_837;
wire r2_420;
assign r2_420 = in[1]? r1_840 : r1_839;
wire r2_421;
assign r2_421 = in[1]? r1_842 : r1_841;
wire r2_422;
assign r2_422 = in[1]? r1_844 : r1_843;
wire r2_423;
assign r2_423 = in[1]? r1_846 : r1_845;
wire r2_424;
assign r2_424 = in[1]? r1_848 : r1_847;
wire r2_425;
assign r2_425 = in[1]? r1_850 : r1_849;
wire r2_426;
assign r2_426 = in[1]? r1_852 : r1_851;
wire r2_427;
assign r2_427 = in[1]? r1_854 : r1_853;
wire r2_428;
assign r2_428 = in[1]? r1_856 : r1_855;
wire r2_429;
assign r2_429 = in[1]? r1_858 : r1_857;
wire r2_430;
assign r2_430 = in[1]? r1_860 : r1_859;
wire r2_431;
assign r2_431 = in[1]? r1_862 : r1_861;
wire r2_432;
assign r2_432 = in[1]? r1_864 : r1_863;
wire r2_433;
assign r2_433 = in[1]? r1_866 : r1_865;
wire r2_434;
assign r2_434 = in[1]? r1_868 : r1_867;
wire r2_435;
assign r2_435 = in[1]? r1_870 : r1_869;
wire r2_436;
assign r2_436 = in[1]? r1_872 : r1_871;
wire r2_437;
assign r2_437 = in[1]? r1_874 : r1_873;
wire r2_438;
assign r2_438 = in[1]? r1_876 : r1_875;
wire r2_439;
assign r2_439 = in[1]? r1_878 : r1_877;
wire r2_440;
assign r2_440 = in[1]? r1_880 : r1_879;
wire r2_441;
assign r2_441 = in[1]? r1_882 : r1_881;
wire r2_442;
assign r2_442 = in[1]? r1_884 : r1_883;
wire r2_443;
assign r2_443 = in[1]? r1_886 : r1_885;
wire r2_444;
assign r2_444 = in[1]? r1_888 : r1_887;
wire r2_445;
assign r2_445 = in[1]? r1_890 : r1_889;
wire r2_446;
assign r2_446 = in[1]? r1_892 : r1_891;
wire r2_447;
assign r2_447 = in[1]? r1_894 : r1_893;
wire r2_448;
assign r2_448 = in[1]? r1_896 : r1_895;
wire r2_449;
assign r2_449 = in[1]? r1_898 : r1_897;
wire r2_450;
assign r2_450 = in[1]? r1_900 : r1_899;
wire r2_451;
assign r2_451 = in[1]? r1_902 : r1_901;
wire r2_452;
assign r2_452 = in[1]? r1_904 : r1_903;
wire r2_453;
assign r2_453 = in[1]? r1_906 : r1_905;
wire r2_454;
assign r2_454 = in[1]? r1_908 : r1_907;
wire r2_455;
assign r2_455 = in[1]? r1_910 : r1_909;
wire r2_456;
assign r2_456 = in[1]? r1_912 : r1_911;
wire r2_457;
assign r2_457 = in[1]? r1_914 : r1_913;
wire r2_458;
assign r2_458 = in[1]? r1_916 : r1_915;
wire r2_459;
assign r2_459 = in[1]? r1_918 : r1_917;
wire r2_460;
assign r2_460 = in[1]? r1_920 : r1_919;
wire r2_461;
assign r2_461 = in[1]? r1_922 : r1_921;
wire r2_462;
assign r2_462 = in[1]? r1_924 : r1_923;
wire r2_463;
assign r2_463 = in[1]? r1_926 : r1_925;
wire r2_464;
assign r2_464 = in[1]? r1_928 : r1_927;
wire r2_465;
assign r2_465 = in[1]? r1_930 : r1_929;
wire r2_466;
assign r2_466 = in[1]? r1_932 : r1_931;
wire r2_467;
assign r2_467 = in[1]? r1_934 : r1_933;
wire r2_468;
assign r2_468 = in[1]? r1_936 : r1_935;
wire r2_469;
assign r2_469 = in[1]? r1_938 : r1_937;
wire r2_470;
assign r2_470 = in[1]? r1_940 : r1_939;
wire r2_471;
assign r2_471 = in[1]? r1_942 : r1_941;
wire r2_472;
assign r2_472 = in[1]? r1_944 : r1_943;
wire r2_473;
assign r2_473 = in[1]? r1_946 : r1_945;
wire r2_474;
assign r2_474 = in[1]? r1_948 : r1_947;
wire r2_475;
assign r2_475 = in[1]? r1_950 : r1_949;
wire r2_476;
assign r2_476 = in[1]? r1_952 : r1_951;
wire r2_477;
assign r2_477 = in[1]? r1_954 : r1_953;
wire r2_478;
assign r2_478 = in[1]? r1_956 : r1_955;
wire r2_479;
assign r2_479 = in[1]? r1_958 : r1_957;
wire r2_480;
assign r2_480 = in[1]? r1_960 : r1_959;
wire r2_481;
assign r2_481 = in[1]? r1_962 : r1_961;
wire r2_482;
assign r2_482 = in[1]? r1_964 : r1_963;
wire r2_483;
assign r2_483 = in[1]? r1_966 : r1_965;
wire r2_484;
assign r2_484 = in[1]? r1_968 : r1_967;
wire r2_485;
assign r2_485 = in[1]? r1_970 : r1_969;
wire r2_486;
assign r2_486 = in[1]? r1_972 : r1_971;
wire r2_487;
assign r2_487 = in[1]? r1_974 : r1_973;
wire r2_488;
assign r2_488 = in[1]? r1_976 : r1_975;
wire r2_489;
assign r2_489 = in[1]? r1_978 : r1_977;
wire r2_490;
assign r2_490 = in[1]? r1_980 : r1_979;
wire r2_491;
assign r2_491 = in[1]? r1_982 : r1_981;
wire r2_492;
assign r2_492 = in[1]? r1_984 : r1_983;
wire r2_493;
assign r2_493 = in[1]? r1_986 : r1_985;
wire r2_494;
assign r2_494 = in[1]? r1_988 : r1_987;
wire r2_495;
assign r2_495 = in[1]? r1_990 : r1_989;
wire r2_496;
assign r2_496 = in[1]? r1_992 : r1_991;
wire r2_497;
assign r2_497 = in[1]? r1_994 : r1_993;
wire r2_498;
assign r2_498 = in[1]? r1_996 : r1_995;
wire r2_499;
assign r2_499 = in[1]? r1_998 : r1_997;
wire r2_500;
assign r2_500 = in[1]? r1_1000 : r1_999;
wire r2_501;
assign r2_501 = in[1]? r1_1002 : r1_1001;
wire r2_502;
assign r2_502 = in[1]? r1_1004 : r1_1003;
wire r2_503;
assign r2_503 = in[1]? r1_1006 : r1_1005;
wire r2_504;
assign r2_504 = in[1]? r1_1008 : r1_1007;
wire r2_505;
assign r2_505 = in[1]? r1_1010 : r1_1009;
wire r2_506;
assign r2_506 = in[1]? r1_1012 : r1_1011;
wire r2_507;
assign r2_507 = in[1]? r1_1014 : r1_1013;
wire r2_508;
assign r2_508 = in[1]? r1_1016 : r1_1015;
wire r2_509;
assign r2_509 = in[1]? r1_1018 : r1_1017;
wire r2_510;
assign r2_510 = in[1]? r1_1020 : r1_1019;
wire r2_511;
assign r2_511 = in[1]? r1_1022 : r1_1021;
wire r2_512;
assign r2_512 = in[1]? r1_1024 : r1_1023;
wire r2_513;
assign r2_513 = in[1]? r1_1026 : r1_1025;
wire r2_514;
assign r2_514 = in[1]? r1_1028 : r1_1027;
wire r2_515;
assign r2_515 = in[1]? r1_1030 : r1_1029;
wire r2_516;
assign r2_516 = in[1]? r1_1032 : r1_1031;
wire r2_517;
assign r2_517 = in[1]? r1_1034 : r1_1033;
wire r2_518;
assign r2_518 = in[1]? r1_1036 : r1_1035;
wire r2_519;
assign r2_519 = in[1]? r1_1038 : r1_1037;
wire r2_520;
assign r2_520 = in[1]? r1_1040 : r1_1039;
wire r2_521;
assign r2_521 = in[1]? r1_1042 : r1_1041;
wire r2_522;
assign r2_522 = in[1]? r1_1044 : r1_1043;
wire r2_523;
assign r2_523 = in[1]? r1_1046 : r1_1045;
wire r2_524;
assign r2_524 = in[1]? r1_1048 : r1_1047;
wire r2_525;
assign r2_525 = in[1]? r1_1050 : r1_1049;
wire r2_526;
assign r2_526 = in[1]? r1_1052 : r1_1051;
wire r2_527;
assign r2_527 = in[1]? r1_1054 : r1_1053;
wire r2_528;
assign r2_528 = in[1]? r1_1056 : r1_1055;
wire r2_529;
assign r2_529 = in[1]? r1_1058 : r1_1057;
wire r2_530;
assign r2_530 = in[1]? r1_1060 : r1_1059;
wire r2_531;
assign r2_531 = in[1]? r1_1062 : r1_1061;
wire r2_532;
assign r2_532 = in[1]? r1_1064 : r1_1063;
wire r2_533;
assign r2_533 = in[1]? r1_1066 : r1_1065;
wire r2_534;
assign r2_534 = in[1]? r1_1068 : r1_1067;
wire r2_535;
assign r2_535 = in[1]? r1_1070 : r1_1069;
wire r2_536;
assign r2_536 = in[1]? r1_1072 : r1_1071;
wire r2_537;
assign r2_537 = in[1]? r1_1074 : r1_1073;
wire r2_538;
assign r2_538 = in[1]? r1_1076 : r1_1075;
wire r2_539;
assign r2_539 = in[1]? r1_1078 : r1_1077;
wire r2_540;
assign r2_540 = in[1]? r1_1080 : r1_1079;
wire r2_541;
assign r2_541 = in[1]? r1_1082 : r1_1081;
wire r2_542;
assign r2_542 = in[1]? r1_1084 : r1_1083;
wire r2_543;
assign r2_543 = in[1]? r1_1086 : r1_1085;
wire r2_544;
assign r2_544 = in[1]? r1_1088 : r1_1087;
wire r2_545;
assign r2_545 = in[1]? r1_1090 : r1_1089;
wire r2_546;
assign r2_546 = in[1]? r1_1092 : r1_1091;
wire r2_547;
assign r2_547 = in[1]? r1_1094 : r1_1093;
wire r2_548;
assign r2_548 = in[1]? r1_1096 : r1_1095;
wire r2_549;
assign r2_549 = in[1]? r1_1098 : r1_1097;
wire r2_550;
assign r2_550 = in[1]? r1_1100 : r1_1099;
wire r2_551;
assign r2_551 = in[1]? r1_1102 : r1_1101;
wire r2_552;
assign r2_552 = in[1]? r1_1104 : r1_1103;
wire r2_553;
assign r2_553 = in[1]? r1_1106 : r1_1105;
wire r2_554;
assign r2_554 = in[1]? r1_1108 : r1_1107;
wire r2_555;
assign r2_555 = in[1]? r1_1110 : r1_1109;
wire r2_556;
assign r2_556 = in[1]? r1_1112 : r1_1111;
wire r2_557;
assign r2_557 = in[1]? r1_1114 : r1_1113;
wire r2_558;
assign r2_558 = in[1]? r1_1116 : r1_1115;
wire r2_559;
assign r2_559 = in[1]? r1_1118 : r1_1117;
wire r2_560;
assign r2_560 = in[1]? r1_1120 : r1_1119;
wire r2_561;
assign r2_561 = in[1]? r1_1122 : r1_1121;
wire r2_562;
assign r2_562 = in[1]? r1_1124 : r1_1123;
wire r2_563;
assign r2_563 = in[1]? r1_1126 : r1_1125;
wire r2_564;
assign r2_564 = in[1]? r1_1128 : r1_1127;
wire r2_565;
assign r2_565 = in[1]? r1_1130 : r1_1129;
wire r2_566;
assign r2_566 = in[1]? r1_1132 : r1_1131;
wire r2_567;
assign r2_567 = in[1]? r1_1134 : r1_1133;
wire r2_568;
assign r2_568 = in[1]? r1_1136 : r1_1135;
wire r2_569;
assign r2_569 = in[1]? r1_1138 : r1_1137;
wire r2_570;
assign r2_570 = in[1]? r1_1140 : r1_1139;
wire r2_571;
assign r2_571 = in[1]? r1_1142 : r1_1141;
wire r2_572;
assign r2_572 = in[1]? r1_1144 : r1_1143;
wire r2_573;
assign r2_573 = in[1]? r1_1146 : r1_1145;
wire r2_574;
assign r2_574 = in[1]? r1_1148 : r1_1147;
wire r2_575;
assign r2_575 = in[1]? r1_1150 : r1_1149;
wire r2_576;
assign r2_576 = in[1]? r1_1152 : r1_1151;
wire r2_577;
assign r2_577 = in[1]? r1_1154 : r1_1153;
wire r2_578;
assign r2_578 = in[1]? r1_1156 : r1_1155;
wire r2_579;
assign r2_579 = in[1]? r1_1158 : r1_1157;
wire r2_580;
assign r2_580 = in[1]? r1_1160 : r1_1159;
wire r2_581;
assign r2_581 = in[1]? r1_1162 : r1_1161;
wire r2_582;
assign r2_582 = in[1]? r1_1164 : r1_1163;
wire r2_583;
assign r2_583 = in[1]? r1_1166 : r1_1165;
wire r2_584;
assign r2_584 = in[1]? r1_1168 : r1_1167;
wire r2_585;
assign r2_585 = in[1]? r1_1170 : r1_1169;
wire r2_586;
assign r2_586 = in[1]? r1_1172 : r1_1171;
wire r2_587;
assign r2_587 = in[1]? r1_1174 : r1_1173;
wire r2_588;
assign r2_588 = in[1]? r1_1176 : r1_1175;
wire r2_589;
assign r2_589 = in[1]? r1_1178 : r1_1177;
wire r2_590;
assign r2_590 = in[1]? r1_1180 : r1_1179;
wire r2_591;
assign r2_591 = in[1]? r1_1182 : r1_1181;
wire r2_592;
assign r2_592 = in[1]? r1_1184 : r1_1183;
wire r2_593;
assign r2_593 = in[1]? r1_1186 : r1_1185;
wire r2_594;
assign r2_594 = in[1]? r1_1188 : r1_1187;
wire r2_595;
assign r2_595 = in[1]? r1_1190 : r1_1189;
wire r2_596;
assign r2_596 = in[1]? r1_1192 : r1_1191;
wire r2_597;
assign r2_597 = in[1]? r1_1194 : r1_1193;
wire r2_598;
assign r2_598 = in[1]? r1_1196 : r1_1195;
wire r2_599;
assign r2_599 = in[1]? r1_1198 : r1_1197;
wire r2_600;
assign r2_600 = in[1]? r1_1200 : r1_1199;
wire r2_601;
assign r2_601 = in[1]? r1_1202 : r1_1201;
wire r2_602;
assign r2_602 = in[1]? r1_1204 : r1_1203;
wire r2_603;
assign r2_603 = in[1]? r1_1206 : r1_1205;
wire r2_604;
assign r2_604 = in[1]? r1_1208 : r1_1207;
wire r2_605;
assign r2_605 = in[1]? r1_1210 : r1_1209;
wire r2_606;
assign r2_606 = in[1]? r1_1212 : r1_1211;
wire r2_607;
assign r2_607 = in[1]? r1_1214 : r1_1213;
wire r2_608;
assign r2_608 = in[1]? r1_1216 : r1_1215;
wire r2_609;
assign r2_609 = in[1]? r1_1218 : r1_1217;
wire r2_610;
assign r2_610 = in[1]? r1_1220 : r1_1219;
wire r2_611;
assign r2_611 = in[1]? r1_1222 : r1_1221;
wire r2_612;
assign r2_612 = in[1]? r1_1224 : r1_1223;
wire r2_613;
assign r2_613 = in[1]? r1_1226 : r1_1225;
wire r2_614;
assign r2_614 = in[1]? r1_1228 : r1_1227;
wire r2_615;
assign r2_615 = in[1]? r1_1230 : r1_1229;
wire r2_616;
assign r2_616 = in[1]? r1_1232 : r1_1231;
wire r2_617;
assign r2_617 = in[1]? r1_1234 : r1_1233;
wire r2_618;
assign r2_618 = in[1]? r1_1236 : r1_1235;
wire r2_619;
assign r2_619 = in[1]? r1_1238 : r1_1237;
wire r2_620;
assign r2_620 = in[1]? r1_1240 : r1_1239;
wire r2_621;
assign r2_621 = in[1]? r1_1242 : r1_1241;
wire r2_622;
assign r2_622 = in[1]? r1_1244 : r1_1243;
wire r2_623;
assign r2_623 = in[1]? r1_1246 : r1_1245;
wire r2_624;
assign r2_624 = in[1]? r1_1248 : r1_1247;
wire r2_625;
assign r2_625 = in[1]? r1_1250 : r1_1249;
wire r2_626;
assign r2_626 = in[1]? r1_1252 : r1_1251;
wire r2_627;
assign r2_627 = in[1]? r1_1254 : r1_1253;
wire r2_628;
assign r2_628 = in[1]? r1_1256 : r1_1255;
wire r2_629;
assign r2_629 = in[1]? r1_1258 : r1_1257;
wire r2_630;
assign r2_630 = in[1]? r1_1260 : r1_1259;
wire r2_631;
assign r2_631 = in[1]? r1_1262 : r1_1261;
wire r2_632;
assign r2_632 = in[1]? r1_1264 : r1_1263;
wire r2_633;
assign r2_633 = in[1]? r1_1266 : r1_1265;
wire r2_634;
assign r2_634 = in[1]? r1_1268 : r1_1267;
wire r2_635;
assign r2_635 = in[1]? r1_1270 : r1_1269;
wire r2_636;
assign r2_636 = in[1]? r1_1272 : r1_1271;
wire r2_637;
assign r2_637 = in[1]? r1_1274 : r1_1273;
wire r2_638;
assign r2_638 = in[1]? r1_1276 : r1_1275;
wire r2_639;
assign r2_639 = in[1]? r1_1278 : r1_1277;
wire r2_640;
assign r2_640 = in[1]? r1_1280 : r1_1279;
wire r2_641;
assign r2_641 = in[1]? r1_1282 : r1_1281;
wire r2_642;
assign r2_642 = in[1]? r1_1284 : r1_1283;
wire r2_643;
assign r2_643 = in[1]? r1_1286 : r1_1285;
wire r2_644;
assign r2_644 = in[1]? r1_1288 : r1_1287;
wire r2_645;
assign r2_645 = in[1]? r1_1290 : r1_1289;
wire r2_646;
assign r2_646 = in[1]? r1_1292 : r1_1291;
wire r2_647;
assign r2_647 = in[1]? r1_1294 : r1_1293;
wire r2_648;
assign r2_648 = in[1]? r1_1296 : r1_1295;
wire r2_649;
assign r2_649 = in[1]? r1_1298 : r1_1297;
wire r2_650;
assign r2_650 = in[1]? r1_1300 : r1_1299;
wire r2_651;
assign r2_651 = in[1]? r1_1302 : r1_1301;
wire r2_652;
assign r2_652 = in[1]? r1_1304 : r1_1303;
wire r2_653;
assign r2_653 = in[1]? r1_1306 : r1_1305;
wire r2_654;
assign r2_654 = in[1]? r1_1308 : r1_1307;
wire r2_655;
assign r2_655 = in[1]? r1_1310 : r1_1309;
wire r2_656;
assign r2_656 = in[1]? r1_1312 : r1_1311;
wire r2_657;
assign r2_657 = in[1]? r1_1314 : r1_1313;
wire r2_658;
assign r2_658 = in[1]? r1_1316 : r1_1315;
wire r2_659;
assign r2_659 = in[1]? r1_1318 : r1_1317;
wire r2_660;
assign r2_660 = in[1]? r1_1320 : r1_1319;
wire r2_661;
assign r2_661 = in[1]? r1_1322 : r1_1321;
wire r2_662;
assign r2_662 = in[1]? r1_1324 : r1_1323;
wire r2_663;
assign r2_663 = in[1]? r1_1326 : r1_1325;
wire r2_664;
assign r2_664 = in[1]? r1_1328 : r1_1327;
wire r2_665;
assign r2_665 = in[1]? r1_1330 : r1_1329;
wire r2_666;
assign r2_666 = in[1]? r1_1332 : r1_1331;
wire r2_667;
assign r2_667 = in[1]? r1_1334 : r1_1333;
wire r2_668;
assign r2_668 = in[1]? r1_1336 : r1_1335;
wire r2_669;
assign r2_669 = in[1]? r1_1338 : r1_1337;
wire r2_670;
assign r2_670 = in[1]? r1_1340 : r1_1339;
wire r2_671;
assign r2_671 = in[1]? r1_1342 : r1_1341;
wire r2_672;
assign r2_672 = in[1]? r1_1344 : r1_1343;
wire r2_673;
assign r2_673 = in[1]? r1_1346 : r1_1345;
wire r2_674;
assign r2_674 = in[1]? r1_1348 : r1_1347;
wire r2_675;
assign r2_675 = in[1]? r1_1350 : r1_1349;
wire r2_676;
assign r2_676 = in[1]? r1_1352 : r1_1351;
wire r2_677;
assign r2_677 = in[1]? r1_1354 : r1_1353;
wire r2_678;
assign r2_678 = in[1]? r1_1356 : r1_1355;
wire r2_679;
assign r2_679 = in[1]? r1_1358 : r1_1357;
wire r2_680;
assign r2_680 = in[1]? r1_1360 : r1_1359;
wire r2_681;
assign r2_681 = in[1]? r1_1362 : r1_1361;
wire r2_682;
assign r2_682 = in[1]? r1_1364 : r1_1363;
wire r2_683;
assign r2_683 = in[1]? r1_1366 : r1_1365;
wire r2_684;
assign r2_684 = in[1]? r1_1368 : r1_1367;
wire r2_685;
assign r2_685 = in[1]? r1_1370 : r1_1369;
wire r2_686;
assign r2_686 = in[1]? r1_1372 : r1_1371;
wire r2_687;
assign r2_687 = in[1]? r1_1374 : r1_1373;
wire r2_688;
assign r2_688 = in[1]? r1_1376 : r1_1375;
wire r2_689;
assign r2_689 = in[1]? r1_1378 : r1_1377;
wire r2_690;
assign r2_690 = in[1]? r1_1380 : r1_1379;
wire r2_691;
assign r2_691 = in[1]? r1_1382 : r1_1381;
wire r2_692;
assign r2_692 = in[1]? r1_1384 : r1_1383;
wire r2_693;
assign r2_693 = in[1]? r1_1386 : r1_1385;
wire r2_694;
assign r2_694 = in[1]? r1_1388 : r1_1387;
wire r2_695;
assign r2_695 = in[1]? r1_1390 : r1_1389;
wire r2_696;
assign r2_696 = in[1]? r1_1392 : r1_1391;
wire r2_697;
assign r2_697 = in[1]? r1_1394 : r1_1393;
wire r2_698;
assign r2_698 = in[1]? r1_1396 : r1_1395;
wire r2_699;
assign r2_699 = in[1]? r1_1398 : r1_1397;
wire r2_700;
assign r2_700 = in[1]? r1_1400 : r1_1399;
wire r2_701;
assign r2_701 = in[1]? r1_1402 : r1_1401;
wire r2_702;
assign r2_702 = in[1]? r1_1404 : r1_1403;
wire r2_703;
assign r2_703 = in[1]? r1_1406 : r1_1405;
wire r2_704;
assign r2_704 = in[1]? r1_1408 : r1_1407;
wire r2_705;
assign r2_705 = in[1]? r1_1410 : r1_1409;
wire r2_706;
assign r2_706 = in[1]? r1_1412 : r1_1411;
wire r2_707;
assign r2_707 = in[1]? r1_1414 : r1_1413;
wire r2_708;
assign r2_708 = in[1]? r1_1416 : r1_1415;
wire r2_709;
assign r2_709 = in[1]? r1_1418 : r1_1417;
wire r2_710;
assign r2_710 = in[1]? r1_1420 : r1_1419;
wire r2_711;
assign r2_711 = in[1]? r1_1422 : r1_1421;
wire r2_712;
assign r2_712 = in[1]? r1_1424 : r1_1423;
wire r2_713;
assign r2_713 = in[1]? r1_1426 : r1_1425;
wire r2_714;
assign r2_714 = in[1]? r1_1428 : r1_1427;
wire r2_715;
assign r2_715 = in[1]? r1_1430 : r1_1429;
wire r2_716;
assign r2_716 = in[1]? r1_1432 : r1_1431;
wire r2_717;
assign r2_717 = in[1]? r1_1434 : r1_1433;
wire r2_718;
assign r2_718 = in[1]? r1_1436 : r1_1435;
wire r2_719;
assign r2_719 = in[1]? r1_1438 : r1_1437;
wire r2_720;
assign r2_720 = in[1]? r1_1440 : r1_1439;
wire r2_721;
assign r2_721 = in[1]? r1_1442 : r1_1441;
wire r2_722;
assign r2_722 = in[1]? r1_1444 : r1_1443;
wire r2_723;
assign r2_723 = in[1]? r1_1446 : r1_1445;
wire r2_724;
assign r2_724 = in[1]? r1_1448 : r1_1447;
wire r2_725;
assign r2_725 = in[1]? r1_1450 : r1_1449;
wire r2_726;
assign r2_726 = in[1]? r1_1452 : r1_1451;
wire r2_727;
assign r2_727 = in[1]? r1_1454 : r1_1453;
wire r2_728;
assign r2_728 = in[1]? r1_1456 : r1_1455;
wire r2_729;
assign r2_729 = in[1]? r1_1458 : r1_1457;
wire r2_730;
assign r2_730 = in[1]? r1_1460 : r1_1459;
wire r2_731;
assign r2_731 = in[1]? r1_1462 : r1_1461;
wire r2_732;
assign r2_732 = in[1]? r1_1464 : r1_1463;
wire r2_733;
assign r2_733 = in[1]? r1_1466 : r1_1465;
wire r2_734;
assign r2_734 = in[1]? r1_1468 : r1_1467;
wire r2_735;
assign r2_735 = in[1]? r1_1470 : r1_1469;
wire r2_736;
assign r2_736 = in[1]? r1_1472 : r1_1471;
wire r2_737;
assign r2_737 = in[1]? r1_1474 : r1_1473;
wire r2_738;
assign r2_738 = in[1]? r1_1476 : r1_1475;
wire r2_739;
assign r2_739 = in[1]? r1_1478 : r1_1477;
wire r2_740;
assign r2_740 = in[1]? r1_1480 : r1_1479;
wire r2_741;
assign r2_741 = in[1]? r1_1482 : r1_1481;
wire r2_742;
assign r2_742 = in[1]? r1_1484 : r1_1483;
wire r2_743;
assign r2_743 = in[1]? r1_1486 : r1_1485;
wire r2_744;
assign r2_744 = in[1]? r1_1488 : r1_1487;
wire r2_745;
assign r2_745 = in[1]? r1_1490 : r1_1489;
wire r2_746;
assign r2_746 = in[1]? r1_1492 : r1_1491;
wire r2_747;
assign r2_747 = in[1]? r1_1494 : r1_1493;
wire r2_748;
assign r2_748 = in[1]? r1_1496 : r1_1495;
wire r2_749;
assign r2_749 = in[1]? r1_1498 : r1_1497;
wire r2_750;
assign r2_750 = in[1]? r1_1500 : r1_1499;
wire r2_751;
assign r2_751 = in[1]? r1_1502 : r1_1501;
wire r2_752;
assign r2_752 = in[1]? r1_1504 : r1_1503;
wire r2_753;
assign r2_753 = in[1]? r1_1506 : r1_1505;
wire r2_754;
assign r2_754 = in[1]? r1_1508 : r1_1507;
wire r2_755;
assign r2_755 = in[1]? r1_1510 : r1_1509;
wire r2_756;
assign r2_756 = in[1]? r1_1512 : r1_1511;
wire r2_757;
assign r2_757 = in[1]? r1_1514 : r1_1513;
wire r2_758;
assign r2_758 = in[1]? r1_1516 : r1_1515;
wire r2_759;
assign r2_759 = in[1]? r1_1518 : r1_1517;
wire r2_760;
assign r2_760 = in[1]? r1_1520 : r1_1519;
wire r2_761;
assign r2_761 = in[1]? r1_1522 : r1_1521;
wire r2_762;
assign r2_762 = in[1]? r1_1524 : r1_1523;
wire r2_763;
assign r2_763 = in[1]? r1_1526 : r1_1525;
wire r2_764;
assign r2_764 = in[1]? r1_1528 : r1_1527;
wire r2_765;
assign r2_765 = in[1]? r1_1530 : r1_1529;
wire r2_766;
assign r2_766 = in[1]? r1_1532 : r1_1531;
wire r2_767;
assign r2_767 = in[1]? r1_1534 : r1_1533;
wire r2_768;
assign r2_768 = in[1]? r1_1536 : r1_1535;
wire r2_769;
assign r2_769 = in[1]? r1_1538 : r1_1537;
wire r2_770;
assign r2_770 = in[1]? r1_1540 : r1_1539;
wire r2_771;
assign r2_771 = in[1]? r1_1542 : r1_1541;
wire r2_772;
assign r2_772 = in[1]? r1_1544 : r1_1543;
wire r2_773;
assign r2_773 = in[1]? r1_1546 : r1_1545;
wire r2_774;
assign r2_774 = in[1]? r1_1548 : r1_1547;
wire r2_775;
assign r2_775 = in[1]? r1_1550 : r1_1549;
wire r2_776;
assign r2_776 = in[1]? r1_1552 : r1_1551;
wire r2_777;
assign r2_777 = in[1]? r1_1554 : r1_1553;
wire r2_778;
assign r2_778 = in[1]? r1_1556 : r1_1555;
wire r2_779;
assign r2_779 = in[1]? r1_1558 : r1_1557;
wire r2_780;
assign r2_780 = in[1]? r1_1560 : r1_1559;
wire r2_781;
assign r2_781 = in[1]? r1_1562 : r1_1561;
wire r2_782;
assign r2_782 = in[1]? r1_1564 : r1_1563;
wire r2_783;
assign r2_783 = in[1]? r1_1566 : r1_1565;
wire r2_784;
assign r2_784 = in[1]? r1_1568 : r1_1567;
wire r2_785;
assign r2_785 = in[1]? r1_1570 : r1_1569;
wire r2_786;
assign r2_786 = in[1]? r1_1572 : r1_1571;
wire r2_787;
assign r2_787 = in[1]? r1_1574 : r1_1573;
wire r2_788;
assign r2_788 = in[1]? r1_1576 : r1_1575;
wire r2_789;
assign r2_789 = in[1]? r1_1578 : r1_1577;
wire r2_790;
assign r2_790 = in[1]? r1_1580 : r1_1579;
wire r2_791;
assign r2_791 = in[1]? r1_1582 : r1_1581;
wire r2_792;
assign r2_792 = in[1]? r1_1584 : r1_1583;
wire r2_793;
assign r2_793 = in[1]? r1_1586 : r1_1585;
wire r2_794;
assign r2_794 = in[1]? r1_1588 : r1_1587;
wire r2_795;
assign r2_795 = in[1]? r1_1590 : r1_1589;
wire r2_796;
assign r2_796 = in[1]? r1_1592 : r1_1591;
wire r2_797;
assign r2_797 = in[1]? r1_1594 : r1_1593;
wire r2_798;
assign r2_798 = in[1]? r1_1596 : r1_1595;
wire r2_799;
assign r2_799 = in[1]? r1_1598 : r1_1597;
wire r2_800;
assign r2_800 = in[1]? r1_1600 : r1_1599;
wire r2_801;
assign r2_801 = in[1]? r1_1602 : r1_1601;
wire r2_802;
assign r2_802 = in[1]? r1_1604 : r1_1603;
wire r2_803;
assign r2_803 = in[1]? r1_1606 : r1_1605;
wire r2_804;
assign r2_804 = in[1]? r1_1608 : r1_1607;
wire r2_805;
assign r2_805 = in[1]? r1_1610 : r1_1609;
wire r2_806;
assign r2_806 = in[1]? r1_1612 : r1_1611;
wire r2_807;
assign r2_807 = in[1]? r1_1614 : r1_1613;
wire r2_808;
assign r2_808 = in[1]? r1_1616 : r1_1615;
wire r2_809;
assign r2_809 = in[1]? r1_1618 : r1_1617;
wire r2_810;
assign r2_810 = in[1]? r1_1620 : r1_1619;
wire r2_811;
assign r2_811 = in[1]? r1_1622 : r1_1621;
wire r2_812;
assign r2_812 = in[1]? r1_1624 : r1_1623;
wire r2_813;
assign r2_813 = in[1]? r1_1626 : r1_1625;
wire r2_814;
assign r2_814 = in[1]? r1_1628 : r1_1627;
wire r2_815;
assign r2_815 = in[1]? r1_1630 : r1_1629;
wire r2_816;
assign r2_816 = in[1]? r1_1632 : r1_1631;
wire r2_817;
assign r2_817 = in[1]? r1_1634 : r1_1633;
wire r2_818;
assign r2_818 = in[1]? r1_1636 : r1_1635;
wire r2_819;
assign r2_819 = in[1]? r1_1638 : r1_1637;
wire r2_820;
assign r2_820 = in[1]? r1_1640 : r1_1639;
wire r2_821;
assign r2_821 = in[1]? r1_1642 : r1_1641;
wire r2_822;
assign r2_822 = in[1]? r1_1644 : r1_1643;
wire r2_823;
assign r2_823 = in[1]? r1_1646 : r1_1645;
wire r2_824;
assign r2_824 = in[1]? r1_1648 : r1_1647;
wire r2_825;
assign r2_825 = in[1]? r1_1650 : r1_1649;
wire r2_826;
assign r2_826 = in[1]? r1_1652 : r1_1651;
wire r2_827;
assign r2_827 = in[1]? r1_1654 : r1_1653;
wire r2_828;
assign r2_828 = in[1]? r1_1656 : r1_1655;
wire r2_829;
assign r2_829 = in[1]? r1_1658 : r1_1657;
wire r2_830;
assign r2_830 = in[1]? r1_1660 : r1_1659;
wire r2_831;
assign r2_831 = in[1]? r1_1662 : r1_1661;
wire r2_832;
assign r2_832 = in[1]? r1_1664 : r1_1663;
wire r2_833;
assign r2_833 = in[1]? r1_1666 : r1_1665;
wire r2_834;
assign r2_834 = in[1]? r1_1668 : r1_1667;
wire r2_835;
assign r2_835 = in[1]? r1_1670 : r1_1669;
wire r2_836;
assign r2_836 = in[1]? r1_1672 : r1_1671;
wire r2_837;
assign r2_837 = in[1]? r1_1674 : r1_1673;
wire r2_838;
assign r2_838 = in[1]? r1_1676 : r1_1675;
wire r2_839;
assign r2_839 = in[1]? r1_1678 : r1_1677;
wire r2_840;
assign r2_840 = in[1]? r1_1680 : r1_1679;
wire r2_841;
assign r2_841 = in[1]? r1_1682 : r1_1681;
wire r2_842;
assign r2_842 = in[1]? r1_1684 : r1_1683;
wire r2_843;
assign r2_843 = in[1]? r1_1686 : r1_1685;
wire r2_844;
assign r2_844 = in[1]? r1_1688 : r1_1687;
wire r2_845;
assign r2_845 = in[1]? r1_1690 : r1_1689;
wire r2_846;
assign r2_846 = in[1]? r1_1692 : r1_1691;
wire r2_847;
assign r2_847 = in[1]? r1_1694 : r1_1693;
wire r2_848;
assign r2_848 = in[1]? r1_1696 : r1_1695;
wire r2_849;
assign r2_849 = in[1]? r1_1698 : r1_1697;
wire r2_850;
assign r2_850 = in[1]? r1_1700 : r1_1699;
wire r2_851;
assign r2_851 = in[1]? r1_1702 : r1_1701;
wire r2_852;
assign r2_852 = in[1]? r1_1704 : r1_1703;
wire r2_853;
assign r2_853 = in[1]? r1_1706 : r1_1705;
wire r2_854;
assign r2_854 = in[1]? r1_1708 : r1_1707;
wire r2_855;
assign r2_855 = in[1]? r1_1710 : r1_1709;
wire r2_856;
assign r2_856 = in[1]? r1_1712 : r1_1711;
wire r2_857;
assign r2_857 = in[1]? r1_1714 : r1_1713;
wire r2_858;
assign r2_858 = in[1]? r1_1716 : r1_1715;
wire r2_859;
assign r2_859 = in[1]? r1_1718 : r1_1717;
wire r2_860;
assign r2_860 = in[1]? r1_1720 : r1_1719;
wire r2_861;
assign r2_861 = in[1]? r1_1722 : r1_1721;
wire r2_862;
assign r2_862 = in[1]? r1_1724 : r1_1723;
wire r2_863;
assign r2_863 = in[1]? r1_1726 : r1_1725;
wire r2_864;
assign r2_864 = in[1]? r1_1728 : r1_1727;
wire r2_865;
assign r2_865 = in[1]? r1_1730 : r1_1729;
wire r2_866;
assign r2_866 = in[1]? r1_1732 : r1_1731;
wire r2_867;
assign r2_867 = in[1]? r1_1734 : r1_1733;
wire r2_868;
assign r2_868 = in[1]? r1_1736 : r1_1735;
wire r2_869;
assign r2_869 = in[1]? r1_1738 : r1_1737;
wire r2_870;
assign r2_870 = in[1]? r1_1740 : r1_1739;
wire r2_871;
assign r2_871 = in[1]? r1_1742 : r1_1741;
wire r2_872;
assign r2_872 = in[1]? r1_1744 : r1_1743;
wire r2_873;
assign r2_873 = in[1]? r1_1746 : r1_1745;
wire r2_874;
assign r2_874 = in[1]? r1_1748 : r1_1747;
wire r2_875;
assign r2_875 = in[1]? r1_1750 : r1_1749;
wire r2_876;
assign r2_876 = in[1]? r1_1752 : r1_1751;
wire r2_877;
assign r2_877 = in[1]? r1_1754 : r1_1753;
wire r2_878;
assign r2_878 = in[1]? r1_1756 : r1_1755;
wire r2_879;
assign r2_879 = in[1]? r1_1758 : r1_1757;
wire r2_880;
assign r2_880 = in[1]? r1_1760 : r1_1759;
wire r2_881;
assign r2_881 = in[1]? r1_1762 : r1_1761;
wire r2_882;
assign r2_882 = in[1]? r1_1764 : r1_1763;
wire r2_883;
assign r2_883 = in[1]? r1_1766 : r1_1765;
wire r2_884;
assign r2_884 = in[1]? r1_1768 : r1_1767;
wire r2_885;
assign r2_885 = in[1]? r1_1770 : r1_1769;
wire r2_886;
assign r2_886 = in[1]? r1_1772 : r1_1771;
wire r2_887;
assign r2_887 = in[1]? r1_1774 : r1_1773;
wire r2_888;
assign r2_888 = in[1]? r1_1776 : r1_1775;
wire r2_889;
assign r2_889 = in[1]? r1_1778 : r1_1777;
wire r2_890;
assign r2_890 = in[1]? r1_1780 : r1_1779;
wire r2_891;
assign r2_891 = in[1]? r1_1782 : r1_1781;
wire r2_892;
assign r2_892 = in[1]? r1_1784 : r1_1783;
wire r2_893;
assign r2_893 = in[1]? r1_1786 : r1_1785;
wire r2_894;
assign r2_894 = in[1]? r1_1788 : r1_1787;
wire r2_895;
assign r2_895 = in[1]? r1_1790 : r1_1789;
wire r2_896;
assign r2_896 = in[1]? r1_1792 : r1_1791;
wire r2_897;
assign r2_897 = in[1]? r1_1794 : r1_1793;
wire r2_898;
assign r2_898 = in[1]? r1_1796 : r1_1795;
wire r2_899;
assign r2_899 = in[1]? r1_1798 : r1_1797;
wire r2_900;
assign r2_900 = in[1]? r1_1800 : r1_1799;
wire r2_901;
assign r2_901 = in[1]? r1_1802 : r1_1801;
wire r2_902;
assign r2_902 = in[1]? r1_1804 : r1_1803;
wire r2_903;
assign r2_903 = in[1]? r1_1806 : r1_1805;
wire r2_904;
assign r2_904 = in[1]? r1_1808 : r1_1807;
wire r2_905;
assign r2_905 = in[1]? r1_1810 : r1_1809;
wire r2_906;
assign r2_906 = in[1]? r1_1812 : r1_1811;
wire r2_907;
assign r2_907 = in[1]? r1_1814 : r1_1813;
wire r2_908;
assign r2_908 = in[1]? r1_1816 : r1_1815;
wire r2_909;
assign r2_909 = in[1]? r1_1818 : r1_1817;
wire r2_910;
assign r2_910 = in[1]? r1_1820 : r1_1819;
wire r2_911;
assign r2_911 = in[1]? r1_1822 : r1_1821;
wire r2_912;
assign r2_912 = in[1]? r1_1824 : r1_1823;
wire r2_913;
assign r2_913 = in[1]? r1_1826 : r1_1825;
wire r2_914;
assign r2_914 = in[1]? r1_1828 : r1_1827;
wire r2_915;
assign r2_915 = in[1]? r1_1830 : r1_1829;
wire r2_916;
assign r2_916 = in[1]? r1_1832 : r1_1831;
wire r2_917;
assign r2_917 = in[1]? r1_1834 : r1_1833;
wire r2_918;
assign r2_918 = in[1]? r1_1836 : r1_1835;
wire r2_919;
assign r2_919 = in[1]? r1_1838 : r1_1837;
wire r2_920;
assign r2_920 = in[1]? r1_1840 : r1_1839;
wire r2_921;
assign r2_921 = in[1]? r1_1842 : r1_1841;
wire r2_922;
assign r2_922 = in[1]? r1_1844 : r1_1843;
wire r2_923;
assign r2_923 = in[1]? r1_1846 : r1_1845;
wire r2_924;
assign r2_924 = in[1]? r1_1848 : r1_1847;
wire r2_925;
assign r2_925 = in[1]? r1_1850 : r1_1849;
wire r2_926;
assign r2_926 = in[1]? r1_1852 : r1_1851;
wire r2_927;
assign r2_927 = in[1]? r1_1854 : r1_1853;
wire r2_928;
assign r2_928 = in[1]? r1_1856 : r1_1855;
wire r2_929;
assign r2_929 = in[1]? r1_1858 : r1_1857;
wire r2_930;
assign r2_930 = in[1]? r1_1860 : r1_1859;
wire r2_931;
assign r2_931 = in[1]? r1_1862 : r1_1861;
wire r2_932;
assign r2_932 = in[1]? r1_1864 : r1_1863;
wire r2_933;
assign r2_933 = in[1]? r1_1866 : r1_1865;
wire r2_934;
assign r2_934 = in[1]? r1_1868 : r1_1867;
wire r2_935;
assign r2_935 = in[1]? r1_1870 : r1_1869;
wire r2_936;
assign r2_936 = in[1]? r1_1872 : r1_1871;
wire r2_937;
assign r2_937 = in[1]? r1_1874 : r1_1873;
wire r2_938;
assign r2_938 = in[1]? r1_1876 : r1_1875;
wire r2_939;
assign r2_939 = in[1]? r1_1878 : r1_1877;
wire r2_940;
assign r2_940 = in[1]? r1_1880 : r1_1879;
wire r2_941;
assign r2_941 = in[1]? r1_1882 : r1_1881;
wire r2_942;
assign r2_942 = in[1]? r1_1884 : r1_1883;
wire r2_943;
assign r2_943 = in[1]? r1_1886 : r1_1885;
wire r2_944;
assign r2_944 = in[1]? r1_1888 : r1_1887;
wire r2_945;
assign r2_945 = in[1]? r1_1890 : r1_1889;
wire r2_946;
assign r2_946 = in[1]? r1_1892 : r1_1891;
wire r2_947;
assign r2_947 = in[1]? r1_1894 : r1_1893;
wire r2_948;
assign r2_948 = in[1]? r1_1896 : r1_1895;
wire r2_949;
assign r2_949 = in[1]? r1_1898 : r1_1897;
wire r2_950;
assign r2_950 = in[1]? r1_1900 : r1_1899;
wire r2_951;
assign r2_951 = in[1]? r1_1902 : r1_1901;
wire r2_952;
assign r2_952 = in[1]? r1_1904 : r1_1903;
wire r2_953;
assign r2_953 = in[1]? r1_1906 : r1_1905;
wire r2_954;
assign r2_954 = in[1]? r1_1908 : r1_1907;
wire r2_955;
assign r2_955 = in[1]? r1_1910 : r1_1909;
wire r2_956;
assign r2_956 = in[1]? r1_1912 : r1_1911;
wire r2_957;
assign r2_957 = in[1]? r1_1914 : r1_1913;
wire r2_958;
assign r2_958 = in[1]? r1_1916 : r1_1915;
wire r2_959;
assign r2_959 = in[1]? r1_1918 : r1_1917;
wire r2_960;
assign r2_960 = in[1]? r1_1920 : r1_1919;
wire r2_961;
assign r2_961 = in[1]? r1_1922 : r1_1921;
wire r2_962;
assign r2_962 = in[1]? r1_1924 : r1_1923;
wire r2_963;
assign r2_963 = in[1]? r1_1926 : r1_1925;
wire r2_964;
assign r2_964 = in[1]? r1_1928 : r1_1927;
wire r2_965;
assign r2_965 = in[1]? r1_1930 : r1_1929;
wire r2_966;
assign r2_966 = in[1]? r1_1932 : r1_1931;
wire r2_967;
assign r2_967 = in[1]? r1_1934 : r1_1933;
wire r2_968;
assign r2_968 = in[1]? r1_1936 : r1_1935;
wire r2_969;
assign r2_969 = in[1]? r1_1938 : r1_1937;
wire r2_970;
assign r2_970 = in[1]? r1_1940 : r1_1939;
wire r2_971;
assign r2_971 = in[1]? r1_1942 : r1_1941;
wire r2_972;
assign r2_972 = in[1]? r1_1944 : r1_1943;
wire r2_973;
assign r2_973 = in[1]? r1_1946 : r1_1945;
wire r2_974;
assign r2_974 = in[1]? r1_1948 : r1_1947;
wire r2_975;
assign r2_975 = in[1]? r1_1950 : r1_1949;
wire r2_976;
assign r2_976 = in[1]? r1_1952 : r1_1951;
wire r2_977;
assign r2_977 = in[1]? r1_1954 : r1_1953;
wire r2_978;
assign r2_978 = in[1]? r1_1956 : r1_1955;
wire r2_979;
assign r2_979 = in[1]? r1_1958 : r1_1957;
wire r2_980;
assign r2_980 = in[1]? r1_1960 : r1_1959;
wire r2_981;
assign r2_981 = in[1]? r1_1962 : r1_1961;
wire r2_982;
assign r2_982 = in[1]? r1_1964 : r1_1963;
wire r2_983;
assign r2_983 = in[1]? r1_1966 : r1_1965;
wire r2_984;
assign r2_984 = in[1]? r1_1968 : r1_1967;
wire r2_985;
assign r2_985 = in[1]? r1_1970 : r1_1969;
wire r2_986;
assign r2_986 = in[1]? r1_1972 : r1_1971;
wire r2_987;
assign r2_987 = in[1]? r1_1974 : r1_1973;
wire r2_988;
assign r2_988 = in[1]? r1_1976 : r1_1975;
wire r2_989;
assign r2_989 = in[1]? r1_1978 : r1_1977;
wire r2_990;
assign r2_990 = in[1]? r1_1980 : r1_1979;
wire r2_991;
assign r2_991 = in[1]? r1_1982 : r1_1981;
wire r2_992;
assign r2_992 = in[1]? r1_1984 : r1_1983;
wire r2_993;
assign r2_993 = in[1]? r1_1986 : r1_1985;
wire r2_994;
assign r2_994 = in[1]? r1_1988 : r1_1987;
wire r2_995;
assign r2_995 = in[1]? r1_1990 : r1_1989;
wire r2_996;
assign r2_996 = in[1]? r1_1992 : r1_1991;
wire r2_997;
assign r2_997 = in[1]? r1_1994 : r1_1993;
wire r2_998;
assign r2_998 = in[1]? r1_1996 : r1_1995;
wire r2_999;
assign r2_999 = in[1]? r1_1998 : r1_1997;
wire r2_1000;
assign r2_1000 = in[1]? r1_2000 : r1_1999;
wire r2_1001;
assign r2_1001 = in[1]? r1_2002 : r1_2001;
wire r2_1002;
assign r2_1002 = in[1]? r1_2004 : r1_2003;
wire r2_1003;
assign r2_1003 = in[1]? r1_2006 : r1_2005;
wire r2_1004;
assign r2_1004 = in[1]? r1_2008 : r1_2007;
wire r2_1005;
assign r2_1005 = in[1]? r1_2010 : r1_2009;
wire r2_1006;
assign r2_1006 = in[1]? r1_2012 : r1_2011;
wire r2_1007;
assign r2_1007 = in[1]? r1_2014 : r1_2013;
wire r2_1008;
assign r2_1008 = in[1]? r1_2016 : r1_2015;
wire r2_1009;
assign r2_1009 = in[1]? r1_2018 : r1_2017;
wire r2_1010;
assign r2_1010 = in[1]? r1_2020 : r1_2019;
wire r2_1011;
assign r2_1011 = in[1]? r1_2022 : r1_2021;
wire r2_1012;
assign r2_1012 = in[1]? r1_2024 : r1_2023;
wire r2_1013;
assign r2_1013 = in[1]? r1_2026 : r1_2025;
wire r2_1014;
assign r2_1014 = in[1]? r1_2028 : r1_2027;
wire r2_1015;
assign r2_1015 = in[1]? r1_2030 : r1_2029;
wire r2_1016;
assign r2_1016 = in[1]? r1_2032 : r1_2031;
wire r2_1017;
assign r2_1017 = in[1]? r1_2034 : r1_2033;
wire r2_1018;
assign r2_1018 = in[1]? r1_2036 : r1_2035;
wire r2_1019;
assign r2_1019 = in[1]? r1_2038 : r1_2037;
wire r2_1020;
assign r2_1020 = in[1]? r1_2040 : r1_2039;
wire r2_1021;
assign r2_1021 = in[1]? r1_2042 : r1_2041;
wire r2_1022;
assign r2_1022 = in[1]? r1_2044 : r1_2043;
wire r2_1023;
assign r2_1023 = in[1]? r1_2046 : r1_2045;
wire r2_1024;
assign r2_1024 = in[1]? r1_2048 : r1_2047;
wire r2_1025;
assign r2_1025 = in[1]? r1_2050 : r1_2049;
wire r2_1026;
assign r2_1026 = in[1]? r1_2052 : r1_2051;
wire r2_1027;
assign r2_1027 = in[1]? r1_2054 : r1_2053;
wire r2_1028;
assign r2_1028 = in[1]? r1_2056 : r1_2055;
wire r2_1029;
assign r2_1029 = in[1]? r1_2058 : r1_2057;
wire r2_1030;
assign r2_1030 = in[1]? r1_2060 : r1_2059;
wire r2_1031;
assign r2_1031 = in[1]? r1_2062 : r1_2061;
wire r2_1032;
assign r2_1032 = in[1]? r1_2064 : r1_2063;
wire r2_1033;
assign r2_1033 = in[1]? r1_2066 : r1_2065;
wire r2_1034;
assign r2_1034 = in[1]? r1_2068 : r1_2067;
wire r2_1035;
assign r2_1035 = in[1]? r1_2070 : r1_2069;
wire r2_1036;
assign r2_1036 = in[1]? r1_2072 : r1_2071;
wire r2_1037;
assign r2_1037 = in[1]? r1_2074 : r1_2073;
wire r2_1038;
assign r2_1038 = in[1]? r1_2076 : r1_2075;
wire r2_1039;
assign r2_1039 = in[1]? r1_2078 : r1_2077;
wire r2_1040;
assign r2_1040 = in[1]? r1_2080 : r1_2079;
wire r2_1041;
assign r2_1041 = in[1]? r1_2082 : r1_2081;
wire r2_1042;
assign r2_1042 = in[1]? r1_2084 : r1_2083;
wire r2_1043;
assign r2_1043 = in[1]? r1_2086 : r1_2085;
wire r2_1044;
assign r2_1044 = in[1]? r1_2088 : r1_2087;
wire r2_1045;
assign r2_1045 = in[1]? r1_2090 : r1_2089;
wire r2_1046;
assign r2_1046 = in[1]? r1_2092 : r1_2091;
wire r2_1047;
assign r2_1047 = in[1]? r1_2094 : r1_2093;
wire r2_1048;
assign r2_1048 = in[1]? r1_2096 : r1_2095;
wire r2_1049;
assign r2_1049 = in[1]? r1_2098 : r1_2097;
wire r2_1050;
assign r2_1050 = in[1]? r1_2100 : r1_2099;
wire r2_1051;
assign r2_1051 = in[1]? r1_2102 : r1_2101;
wire r2_1052;
assign r2_1052 = in[1]? r1_2104 : r1_2103;
wire r2_1053;
assign r2_1053 = in[1]? r1_2106 : r1_2105;
wire r2_1054;
assign r2_1054 = in[1]? r1_2108 : r1_2107;
wire r2_1055;
assign r2_1055 = in[1]? r1_2110 : r1_2109;
wire r2_1056;
assign r2_1056 = in[1]? r1_2112 : r1_2111;
wire r2_1057;
assign r2_1057 = in[1]? r1_2114 : r1_2113;
wire r2_1058;
assign r2_1058 = in[1]? r1_2116 : r1_2115;
wire r2_1059;
assign r2_1059 = in[1]? r1_2118 : r1_2117;
wire r2_1060;
assign r2_1060 = in[1]? r1_2120 : r1_2119;
wire r2_1061;
assign r2_1061 = in[1]? r1_2122 : r1_2121;
wire r2_1062;
assign r2_1062 = in[1]? r1_2124 : r1_2123;
wire r2_1063;
assign r2_1063 = in[1]? r1_2126 : r1_2125;
wire r2_1064;
assign r2_1064 = in[1]? r1_2128 : r1_2127;
wire r2_1065;
assign r2_1065 = in[1]? r1_2130 : r1_2129;
wire r2_1066;
assign r2_1066 = in[1]? r1_2132 : r1_2131;
wire r2_1067;
assign r2_1067 = in[1]? r1_2134 : r1_2133;
wire r2_1068;
assign r2_1068 = in[1]? r1_2136 : r1_2135;
wire r2_1069;
assign r2_1069 = in[1]? r1_2138 : r1_2137;
wire r2_1070;
assign r2_1070 = in[1]? r1_2140 : r1_2139;
wire r2_1071;
assign r2_1071 = in[1]? r1_2142 : r1_2141;
wire r2_1072;
assign r2_1072 = in[1]? r1_2144 : r1_2143;
wire r2_1073;
assign r2_1073 = in[1]? r1_2146 : r1_2145;
wire r2_1074;
assign r2_1074 = in[1]? r1_2148 : r1_2147;
wire r2_1075;
assign r2_1075 = in[1]? r1_2150 : r1_2149;
wire r2_1076;
assign r2_1076 = in[1]? r1_2152 : r1_2151;
wire r2_1077;
assign r2_1077 = in[1]? r1_2154 : r1_2153;
wire r2_1078;
assign r2_1078 = in[1]? r1_2156 : r1_2155;
wire r2_1079;
assign r2_1079 = in[1]? r1_2158 : r1_2157;
wire r2_1080;
assign r2_1080 = in[1]? r1_2160 : r1_2159;
wire r2_1081;
assign r2_1081 = in[1]? r1_2162 : r1_2161;
wire r2_1082;
assign r2_1082 = in[1]? r1_2164 : r1_2163;
wire r2_1083;
assign r2_1083 = in[1]? r1_2166 : r1_2165;
wire r2_1084;
assign r2_1084 = in[1]? r1_2168 : r1_2167;
wire r2_1085;
assign r2_1085 = in[1]? r1_2170 : r1_2169;
wire r2_1086;
assign r2_1086 = in[1]? r1_2172 : r1_2171;
wire r2_1087;
assign r2_1087 = in[1]? r1_2174 : r1_2173;
wire r2_1088;
assign r2_1088 = in[1]? r1_2176 : r1_2175;
wire r2_1089;
assign r2_1089 = in[1]? r1_2178 : r1_2177;
wire r2_1090;
assign r2_1090 = in[1]? r1_2180 : r1_2179;
wire r2_1091;
assign r2_1091 = in[1]? r1_2182 : r1_2181;
wire r2_1092;
assign r2_1092 = in[1]? r1_2184 : r1_2183;
wire r2_1093;
assign r2_1093 = in[1]? r1_2186 : r1_2185;
wire r2_1094;
assign r2_1094 = in[1]? r1_2188 : r1_2187;
wire r2_1095;
assign r2_1095 = in[1]? r1_2190 : r1_2189;
wire r2_1096;
assign r2_1096 = in[1]? r1_2192 : r1_2191;
wire r2_1097;
assign r2_1097 = in[1]? r1_2194 : r1_2193;
wire r2_1098;
assign r2_1098 = in[1]? r1_2196 : r1_2195;
wire r2_1099;
assign r2_1099 = in[1]? r1_2198 : r1_2197;
wire r2_1100;
assign r2_1100 = in[1]? r1_2200 : r1_2199;
wire r2_1101;
assign r2_1101 = in[1]? r1_2202 : r1_2201;
wire r2_1102;
assign r2_1102 = in[1]? r1_2204 : r1_2203;
wire r2_1103;
assign r2_1103 = in[1]? r1_2206 : r1_2205;
wire r2_1104;
assign r2_1104 = in[1]? r1_2208 : r1_2207;
wire r2_1105;
assign r2_1105 = in[1]? r1_2210 : r1_2209;
wire r2_1106;
assign r2_1106 = in[1]? r1_2212 : r1_2211;
wire r2_1107;
assign r2_1107 = in[1]? r1_2214 : r1_2213;
wire r2_1108;
assign r2_1108 = in[1]? r1_2216 : r1_2215;
wire r2_1109;
assign r2_1109 = in[1]? r1_2218 : r1_2217;
wire r2_1110;
assign r2_1110 = in[1]? r1_2220 : r1_2219;
wire r2_1111;
assign r2_1111 = in[1]? r1_2222 : r1_2221;
wire r2_1112;
assign r2_1112 = in[1]? r1_2224 : r1_2223;
wire r2_1113;
assign r2_1113 = in[1]? r1_2226 : r1_2225;
wire r2_1114;
assign r2_1114 = in[1]? r1_2228 : r1_2227;
wire r2_1115;
assign r2_1115 = in[1]? r1_2230 : r1_2229;
wire r2_1116;
assign r2_1116 = in[1]? r1_2232 : r1_2231;
wire r2_1117;
assign r2_1117 = in[1]? r1_2234 : r1_2233;
wire r2_1118;
assign r2_1118 = in[1]? r1_2236 : r1_2235;
wire r2_1119;
assign r2_1119 = in[1]? r1_2238 : r1_2237;
wire r2_1120;
assign r2_1120 = in[1]? r1_2240 : r1_2239;
wire r2_1121;
assign r2_1121 = in[1]? r1_2242 : r1_2241;
wire r2_1122;
assign r2_1122 = in[1]? r1_2244 : r1_2243;
wire r2_1123;
assign r2_1123 = in[1]? r1_2246 : r1_2245;
wire r2_1124;
assign r2_1124 = in[1]? r1_2248 : r1_2247;
wire r2_1125;
assign r2_1125 = in[1]? r1_2250 : r1_2249;
wire r2_1126;
assign r2_1126 = in[1]? r1_2252 : r1_2251;
wire r2_1127;
assign r2_1127 = in[1]? r1_2254 : r1_2253;
wire r2_1128;
assign r2_1128 = in[1]? r1_2256 : r1_2255;
wire r2_1129;
assign r2_1129 = in[1]? r1_2258 : r1_2257;
wire r2_1130;
assign r2_1130 = in[1]? r1_2260 : r1_2259;
wire r2_1131;
assign r2_1131 = in[1]? r1_2262 : r1_2261;
wire r2_1132;
assign r2_1132 = in[1]? r1_2264 : r1_2263;
wire r2_1133;
assign r2_1133 = in[1]? r1_2266 : r1_2265;
wire r2_1134;
assign r2_1134 = in[1]? r1_2268 : r1_2267;
wire r2_1135;
assign r2_1135 = in[1]? r1_2270 : r1_2269;
wire r2_1136;
assign r2_1136 = in[1]? r1_2272 : r1_2271;
wire r2_1137;
assign r2_1137 = in[1]? r1_2274 : r1_2273;
wire r2_1138;
assign r2_1138 = in[1]? r1_2276 : r1_2275;
wire r2_1139;
assign r2_1139 = in[1]? r1_2278 : r1_2277;
wire r2_1140;
assign r2_1140 = in[1]? r1_2280 : r1_2279;
wire r2_1141;
assign r2_1141 = in[1]? r1_2282 : r1_2281;
wire r2_1142;
assign r2_1142 = in[1]? r1_2284 : r1_2283;
wire r2_1143;
assign r2_1143 = in[1]? r1_2286 : r1_2285;
wire r2_1144;
assign r2_1144 = in[1]? r1_2288 : r1_2287;
wire r2_1145;
assign r2_1145 = in[1]? r1_2290 : r1_2289;
wire r2_1146;
assign r2_1146 = in[1]? r1_2292 : r1_2291;
wire r2_1147;
assign r2_1147 = in[1]? r1_2294 : r1_2293;
wire r2_1148;
assign r2_1148 = in[1]? r1_2296 : r1_2295;
wire r2_1149;
assign r2_1149 = in[1]? r1_2298 : r1_2297;
wire r2_1150;
assign r2_1150 = in[1]? r1_2300 : r1_2299;
wire r2_1151;
assign r2_1151 = in[1]? r1_2302 : r1_2301;
wire r2_1152;
assign r2_1152 = in[1]? r1_2304 : r1_2303;
wire r2_1153;
assign r2_1153 = in[1]? r1_2306 : r1_2305;
wire r2_1154;
assign r2_1154 = in[1]? r1_2308 : r1_2307;
wire r2_1155;
assign r2_1155 = in[1]? r1_2310 : r1_2309;
wire r2_1156;
assign r2_1156 = in[1]? r1_2312 : r1_2311;
wire r2_1157;
assign r2_1157 = in[1]? r1_2314 : r1_2313;
wire r2_1158;
assign r2_1158 = in[1]? r1_2316 : r1_2315;
wire r2_1159;
assign r2_1159 = in[1]? r1_2318 : r1_2317;
wire r2_1160;
assign r2_1160 = in[1]? r1_2320 : r1_2319;
wire r2_1161;
assign r2_1161 = in[1]? r1_2322 : r1_2321;
wire r2_1162;
assign r2_1162 = in[1]? r1_2324 : r1_2323;
wire r2_1163;
assign r2_1163 = in[1]? r1_2326 : r1_2325;
wire r2_1164;
assign r2_1164 = in[1]? r1_2328 : r1_2327;
wire r2_1165;
assign r2_1165 = in[1]? r1_2330 : r1_2329;
wire r2_1166;
assign r2_1166 = in[1]? r1_2332 : r1_2331;
wire r2_1167;
assign r2_1167 = in[1]? r1_2334 : r1_2333;
wire r2_1168;
assign r2_1168 = in[1]? r1_2336 : r1_2335;
wire r2_1169;
assign r2_1169 = in[1]? r1_2338 : r1_2337;
wire r2_1170;
assign r2_1170 = in[1]? r1_2340 : r1_2339;
wire r2_1171;
assign r2_1171 = in[1]? r1_2342 : r1_2341;
wire r2_1172;
assign r2_1172 = in[1]? r1_2344 : r1_2343;
wire r2_1173;
assign r2_1173 = in[1]? r1_2346 : r1_2345;
wire r2_1174;
assign r2_1174 = in[1]? r1_2348 : r1_2347;
wire r2_1175;
assign r2_1175 = in[1]? r1_2350 : r1_2349;
wire r2_1176;
assign r2_1176 = in[1]? r1_2352 : r1_2351;
wire r2_1177;
assign r2_1177 = in[1]? r1_2354 : r1_2353;
wire r2_1178;
assign r2_1178 = in[1]? r1_2356 : r1_2355;
wire r2_1179;
assign r2_1179 = in[1]? r1_2358 : r1_2357;
wire r2_1180;
assign r2_1180 = in[1]? r1_2360 : r1_2359;
wire r2_1181;
assign r2_1181 = in[1]? r1_2362 : r1_2361;
wire r2_1182;
assign r2_1182 = in[1]? r1_2364 : r1_2363;
wire r2_1183;
assign r2_1183 = in[1]? r1_2366 : r1_2365;
wire r2_1184;
assign r2_1184 = in[1]? r1_2368 : r1_2367;
wire r2_1185;
assign r2_1185 = in[1]? r1_2370 : r1_2369;
wire r2_1186;
assign r2_1186 = in[1]? r1_2372 : r1_2371;
wire r2_1187;
assign r2_1187 = in[1]? r1_2374 : r1_2373;
wire r2_1188;
assign r2_1188 = in[1]? r1_2376 : r1_2375;
wire r2_1189;
assign r2_1189 = in[1]? r1_2378 : r1_2377;
wire r2_1190;
assign r2_1190 = in[1]? r1_2380 : r1_2379;
wire r2_1191;
assign r2_1191 = in[1]? r1_2382 : r1_2381;
wire r2_1192;
assign r2_1192 = in[1]? r1_2384 : r1_2383;
wire r2_1193;
assign r2_1193 = in[1]? r1_2386 : r1_2385;
wire r2_1194;
assign r2_1194 = in[1]? r1_2388 : r1_2387;
wire r2_1195;
assign r2_1195 = in[1]? r1_2390 : r1_2389;
wire r2_1196;
assign r2_1196 = in[1]? r1_2392 : r1_2391;
wire r2_1197;
assign r2_1197 = in[1]? r1_2394 : r1_2393;
wire r2_1198;
assign r2_1198 = in[1]? r1_2396 : r1_2395;
wire r2_1199;
assign r2_1199 = in[1]? r1_2398 : r1_2397;
wire r2_1200;
assign r2_1200 = in[1]? r1_2400 : r1_2399;
wire r2_1201;
assign r2_1201 = in[1]? r1_2402 : r1_2401;
wire r2_1202;
assign r2_1202 = in[1]? r1_2404 : r1_2403;
wire r2_1203;
assign r2_1203 = in[1]? r1_2406 : r1_2405;
wire r2_1204;
assign r2_1204 = in[1]? r1_2408 : r1_2407;
wire r2_1205;
assign r2_1205 = in[1]? r1_2410 : r1_2409;
wire r2_1206;
assign r2_1206 = in[1]? r1_2412 : r1_2411;
wire r2_1207;
assign r2_1207 = in[1]? r1_2414 : r1_2413;
wire r2_1208;
assign r2_1208 = in[1]? r1_2416 : r1_2415;
wire r2_1209;
assign r2_1209 = in[1]? r1_2418 : r1_2417;
wire r2_1210;
assign r2_1210 = in[1]? r1_2420 : r1_2419;
wire r2_1211;
assign r2_1211 = in[1]? r1_2422 : r1_2421;
wire r2_1212;
assign r2_1212 = in[1]? r1_2424 : r1_2423;
wire r2_1213;
assign r2_1213 = in[1]? r1_2426 : r1_2425;
wire r2_1214;
assign r2_1214 = in[1]? r1_2428 : r1_2427;
wire r2_1215;
assign r2_1215 = in[1]? r1_2430 : r1_2429;
wire r2_1216;
assign r2_1216 = in[1]? r1_2432 : r1_2431;
wire r2_1217;
assign r2_1217 = in[1]? r1_2434 : r1_2433;
wire r2_1218;
assign r2_1218 = in[1]? r1_2436 : r1_2435;
wire r2_1219;
assign r2_1219 = in[1]? r1_2438 : r1_2437;
wire r2_1220;
assign r2_1220 = in[1]? r1_2440 : r1_2439;
wire r2_1221;
assign r2_1221 = in[1]? r1_2442 : r1_2441;
wire r2_1222;
assign r2_1222 = in[1]? r1_2444 : r1_2443;
wire r2_1223;
assign r2_1223 = in[1]? r1_2446 : r1_2445;
wire r2_1224;
assign r2_1224 = in[1]? r1_2448 : r1_2447;
wire r2_1225;
assign r2_1225 = in[1]? r1_2450 : r1_2449;
wire r2_1226;
assign r2_1226 = in[1]? r1_2452 : r1_2451;
wire r2_1227;
assign r2_1227 = in[1]? r1_2454 : r1_2453;
wire r2_1228;
assign r2_1228 = in[1]? r1_2456 : r1_2455;
wire r2_1229;
assign r2_1229 = in[1]? r1_2458 : r1_2457;
wire r2_1230;
assign r2_1230 = in[1]? r1_2460 : r1_2459;
wire r2_1231;
assign r2_1231 = in[1]? r1_2462 : r1_2461;
wire r2_1232;
assign r2_1232 = in[1]? r1_2464 : r1_2463;
wire r2_1233;
assign r2_1233 = in[1]? r1_2466 : r1_2465;
wire r2_1234;
assign r2_1234 = in[1]? r1_2468 : r1_2467;
wire r2_1235;
assign r2_1235 = in[1]? r1_2470 : r1_2469;
wire r2_1236;
assign r2_1236 = in[1]? r1_2472 : r1_2471;
wire r2_1237;
assign r2_1237 = in[1]? r1_2474 : r1_2473;
wire r2_1238;
assign r2_1238 = in[1]? r1_2476 : r1_2475;
wire r2_1239;
assign r2_1239 = in[1]? r1_2478 : r1_2477;
wire r2_1240;
assign r2_1240 = in[1]? r1_2480 : r1_2479;
wire r2_1241;
assign r2_1241 = in[1]? r1_2482 : r1_2481;
wire r2_1242;
assign r2_1242 = in[1]? r1_2484 : r1_2483;
wire r2_1243;
assign r2_1243 = in[1]? r1_2486 : r1_2485;
wire r2_1244;
assign r2_1244 = in[1]? r1_2488 : r1_2487;
wire r2_1245;
assign r2_1245 = in[1]? r1_2490 : r1_2489;
wire r2_1246;
assign r2_1246 = in[1]? r1_2492 : r1_2491;
wire r2_1247;
assign r2_1247 = in[1]? r1_2494 : r1_2493;
wire r2_1248;
assign r2_1248 = in[1]? r1_2496 : r1_2495;
wire r2_1249;
assign r2_1249 = in[1]? r1_2498 : r1_2497;
wire r2_1250;
assign r2_1250 = in[1]? r1_2500 : r1_2499;
wire r2_1251;
assign r2_1251 = in[1]? r1_2502 : r1_2501;
wire r2_1252;
assign r2_1252 = in[1]? r1_2504 : r1_2503;
wire r2_1253;
assign r2_1253 = in[1]? r1_2506 : r1_2505;
wire r2_1254;
assign r2_1254 = in[1]? r1_2508 : r1_2507;
wire r2_1255;
assign r2_1255 = in[1]? r1_2510 : r1_2509;
wire r2_1256;
assign r2_1256 = in[1]? r1_2512 : r1_2511;
wire r2_1257;
assign r2_1257 = in[1]? r1_2514 : r1_2513;
wire r2_1258;
assign r2_1258 = in[1]? r1_2516 : r1_2515;
wire r2_1259;
assign r2_1259 = in[1]? r1_2518 : r1_2517;
wire r2_1260;
assign r2_1260 = in[1]? r1_2520 : r1_2519;
wire r2_1261;
assign r2_1261 = in[1]? r1_2522 : r1_2521;
wire r2_1262;
assign r2_1262 = in[1]? r1_2524 : r1_2523;
wire r2_1263;
assign r2_1263 = in[1]? r1_2526 : r1_2525;
wire r2_1264;
assign r2_1264 = in[1]? r1_2528 : r1_2527;
wire r2_1265;
assign r2_1265 = in[1]? r1_2530 : r1_2529;
wire r2_1266;
assign r2_1266 = in[1]? r1_2532 : r1_2531;
wire r2_1267;
assign r2_1267 = in[1]? r1_2534 : r1_2533;
wire r2_1268;
assign r2_1268 = in[1]? r1_2536 : r1_2535;
wire r2_1269;
assign r2_1269 = in[1]? r1_2538 : r1_2537;
wire r2_1270;
assign r2_1270 = in[1]? r1_2540 : r1_2539;
wire r2_1271;
assign r2_1271 = in[1]? r1_2542 : r1_2541;
wire r2_1272;
assign r2_1272 = in[1]? r1_2544 : r1_2543;
wire r2_1273;
assign r2_1273 = in[1]? r1_2546 : r1_2545;
wire r2_1274;
assign r2_1274 = in[1]? r1_2548 : r1_2547;
wire r2_1275;
assign r2_1275 = in[1]? r1_2550 : r1_2549;
wire r2_1276;
assign r2_1276 = in[1]? r1_2552 : r1_2551;
wire r2_1277;
assign r2_1277 = in[1]? r1_2554 : r1_2553;
wire r2_1278;
assign r2_1278 = in[1]? r1_2556 : r1_2555;
wire r2_1279;
assign r2_1279 = in[1]? r1_2558 : r1_2557;
wire r2_1280;
assign r2_1280 = in[1]? r1_2560 : r1_2559;
wire r2_1281;
assign r2_1281 = in[1]? r1_2562 : r1_2561;
wire r2_1282;
assign r2_1282 = in[1]? r1_2564 : r1_2563;
wire r2_1283;
assign r2_1283 = in[1]? r1_2566 : r1_2565;
wire r2_1284;
assign r2_1284 = in[1]? r1_2568 : r1_2567;
wire r2_1285;
assign r2_1285 = in[1]? r1_2570 : r1_2569;
wire r2_1286;
assign r2_1286 = in[1]? r1_2572 : r1_2571;
wire r2_1287;
assign r2_1287 = in[1]? r1_2574 : r1_2573;
wire r2_1288;
assign r2_1288 = in[1]? r1_2576 : r1_2575;
wire r2_1289;
assign r2_1289 = in[1]? r1_2578 : r1_2577;
wire r2_1290;
assign r2_1290 = in[1]? r1_2580 : r1_2579;
wire r2_1291;
assign r2_1291 = in[1]? r1_2582 : r1_2581;
wire r2_1292;
assign r2_1292 = in[1]? r1_2584 : r1_2583;
wire r2_1293;
assign r2_1293 = in[1]? r1_2586 : r1_2585;
wire r2_1294;
assign r2_1294 = in[1]? r1_2588 : r1_2587;
wire r2_1295;
assign r2_1295 = in[1]? r1_2590 : r1_2589;
wire r2_1296;
assign r2_1296 = in[1]? r1_2592 : r1_2591;
wire r2_1297;
assign r2_1297 = in[1]? r1_2594 : r1_2593;
wire r2_1298;
assign r2_1298 = in[1]? r1_2596 : r1_2595;
wire r2_1299;
assign r2_1299 = in[1]? r1_2598 : r1_2597;
wire r2_1300;
assign r2_1300 = in[1]? r1_2600 : r1_2599;
wire r2_1301;
assign r2_1301 = in[1]? r1_2602 : r1_2601;
wire r2_1302;
assign r2_1302 = in[1]? r1_2604 : r1_2603;
wire r2_1303;
assign r2_1303 = in[1]? r1_2606 : r1_2605;
wire r2_1304;
assign r2_1304 = in[1]? r1_2608 : r1_2607;
wire r2_1305;
assign r2_1305 = in[1]? r1_2610 : r1_2609;
wire r2_1306;
assign r2_1306 = in[1]? r1_2612 : r1_2611;
wire r2_1307;
assign r2_1307 = in[1]? r1_2614 : r1_2613;
wire r2_1308;
assign r2_1308 = in[1]? r1_2616 : r1_2615;
wire r2_1309;
assign r2_1309 = in[1]? r1_2618 : r1_2617;
wire r2_1310;
assign r2_1310 = in[1]? r1_2620 : r1_2619;
wire r2_1311;
assign r2_1311 = in[1]? r1_2622 : r1_2621;
wire r2_1312;
assign r2_1312 = in[1]? r1_2624 : r1_2623;
wire r2_1313;
assign r2_1313 = in[1]? r1_2626 : r1_2625;
wire r2_1314;
assign r2_1314 = in[1]? r1_2628 : r1_2627;
wire r2_1315;
assign r2_1315 = in[1]? r1_2630 : r1_2629;
wire r2_1316;
assign r2_1316 = in[1]? r1_2632 : r1_2631;
wire r2_1317;
assign r2_1317 = in[1]? r1_2634 : r1_2633;
wire r2_1318;
assign r2_1318 = in[1]? r1_2636 : r1_2635;
wire r2_1319;
assign r2_1319 = in[1]? r1_2638 : r1_2637;
wire r2_1320;
assign r2_1320 = in[1]? r1_2640 : r1_2639;
wire r2_1321;
assign r2_1321 = in[1]? r1_2642 : r1_2641;
wire r2_1322;
assign r2_1322 = in[1]? r1_2644 : r1_2643;
wire r2_1323;
assign r2_1323 = in[1]? r1_2646 : r1_2645;
wire r2_1324;
assign r2_1324 = in[1]? r1_2648 : r1_2647;
wire r2_1325;
assign r2_1325 = in[1]? r1_2650 : r1_2649;
wire r2_1326;
assign r2_1326 = in[1]? r1_2652 : r1_2651;
wire r2_1327;
assign r2_1327 = in[1]? r1_2654 : r1_2653;
wire r2_1328;
assign r2_1328 = in[1]? r1_2656 : r1_2655;
wire r2_1329;
assign r2_1329 = in[1]? r1_2658 : r1_2657;
wire r2_1330;
assign r2_1330 = in[1]? r1_2660 : r1_2659;
wire r2_1331;
assign r2_1331 = in[1]? r1_2662 : r1_2661;
wire r2_1332;
assign r2_1332 = in[1]? r1_2664 : r1_2663;
wire r2_1333;
assign r2_1333 = in[1]? r1_2666 : r1_2665;
wire r2_1334;
assign r2_1334 = in[1]? r1_2668 : r1_2667;
wire r2_1335;
assign r2_1335 = in[1]? r1_2670 : r1_2669;
wire r2_1336;
assign r2_1336 = in[1]? r1_2672 : r1_2671;
wire r2_1337;
assign r2_1337 = in[1]? r1_2674 : r1_2673;
wire r2_1338;
assign r2_1338 = in[1]? r1_2676 : r1_2675;
wire r2_1339;
assign r2_1339 = in[1]? r1_2678 : r1_2677;
wire r2_1340;
assign r2_1340 = in[1]? r1_2680 : r1_2679;
wire r2_1341;
assign r2_1341 = in[1]? r1_2682 : r1_2681;
wire r2_1342;
assign r2_1342 = in[1]? r1_2684 : r1_2683;
wire r2_1343;
assign r2_1343 = in[1]? r1_2686 : r1_2685;
wire r2_1344;
assign r2_1344 = in[1]? r1_2688 : r1_2687;
wire r2_1345;
assign r2_1345 = in[1]? r1_2690 : r1_2689;
wire r2_1346;
assign r2_1346 = in[1]? r1_2692 : r1_2691;
wire r2_1347;
assign r2_1347 = in[1]? r1_2694 : r1_2693;
wire r2_1348;
assign r2_1348 = in[1]? r1_2696 : r1_2695;
wire r2_1349;
assign r2_1349 = in[1]? r1_2698 : r1_2697;
wire r2_1350;
assign r2_1350 = in[1]? r1_2700 : r1_2699;
wire r2_1351;
assign r2_1351 = in[1]? r1_2702 : r1_2701;
wire r2_1352;
assign r2_1352 = in[1]? r1_2704 : r1_2703;
wire r2_1353;
assign r2_1353 = in[1]? r1_2706 : r1_2705;
wire r2_1354;
assign r2_1354 = in[1]? r1_2708 : r1_2707;
wire r2_1355;
assign r2_1355 = in[1]? r1_2710 : r1_2709;
wire r2_1356;
assign r2_1356 = in[1]? r1_2712 : r1_2711;
wire r2_1357;
assign r2_1357 = in[1]? r1_2714 : r1_2713;
wire r2_1358;
assign r2_1358 = in[1]? r1_2716 : r1_2715;
wire r2_1359;
assign r2_1359 = in[1]? r1_2718 : r1_2717;
wire r2_1360;
assign r2_1360 = in[1]? r1_2720 : r1_2719;
wire r2_1361;
assign r2_1361 = in[1]? r1_2722 : r1_2721;
wire r2_1362;
assign r2_1362 = in[1]? r1_2724 : r1_2723;
wire r2_1363;
assign r2_1363 = in[1]? r1_2726 : r1_2725;
wire r2_1364;
assign r2_1364 = in[1]? r1_2728 : r1_2727;
wire r2_1365;
assign r2_1365 = in[1]? r1_2730 : r1_2729;
wire r2_1366;
assign r2_1366 = in[1]? r1_2732 : r1_2731;
wire r2_1367;
assign r2_1367 = in[1]? r1_2734 : r1_2733;
wire r2_1368;
assign r2_1368 = in[1]? r1_2736 : r1_2735;
wire r2_1369;
assign r2_1369 = in[1]? r1_2738 : r1_2737;
wire r2_1370;
assign r2_1370 = in[1]? r1_2740 : r1_2739;
wire r2_1371;
assign r2_1371 = in[1]? r1_2742 : r1_2741;
wire r2_1372;
assign r2_1372 = in[1]? r1_2744 : r1_2743;
wire r2_1373;
assign r2_1373 = in[1]? r1_2746 : r1_2745;
wire r2_1374;
assign r2_1374 = in[1]? r1_2748 : r1_2747;
wire r2_1375;
assign r2_1375 = in[1]? r1_2750 : r1_2749;
wire r2_1376;
assign r2_1376 = in[1]? r1_2752 : r1_2751;
wire r2_1377;
assign r2_1377 = in[1]? r1_2754 : r1_2753;
wire r2_1378;
assign r2_1378 = in[1]? r1_2756 : r1_2755;
wire r2_1379;
assign r2_1379 = in[1]? r1_2758 : r1_2757;
wire r2_1380;
assign r2_1380 = in[1]? r1_2760 : r1_2759;
wire r2_1381;
assign r2_1381 = in[1]? r1_2762 : r1_2761;
wire r2_1382;
assign r2_1382 = in[1]? r1_2764 : r1_2763;
wire r2_1383;
assign r2_1383 = in[1]? r1_2766 : r1_2765;
wire r2_1384;
assign r2_1384 = in[1]? r1_2768 : r1_2767;
wire r2_1385;
assign r2_1385 = in[1]? r1_2770 : r1_2769;
wire r2_1386;
assign r2_1386 = in[1]? r1_2772 : r1_2771;
wire r2_1387;
assign r2_1387 = in[1]? r1_2774 : r1_2773;
wire r2_1388;
assign r2_1388 = in[1]? r1_2776 : r1_2775;
wire r2_1389;
assign r2_1389 = in[1]? r1_2778 : r1_2777;
wire r2_1390;
assign r2_1390 = in[1]? r1_2780 : r1_2779;
wire r2_1391;
assign r2_1391 = in[1]? r1_2782 : r1_2781;
wire r2_1392;
assign r2_1392 = in[1]? r1_2784 : r1_2783;
wire r2_1393;
assign r2_1393 = in[1]? r1_2786 : r1_2785;
wire r2_1394;
assign r2_1394 = in[1]? r1_2788 : r1_2787;
wire r2_1395;
assign r2_1395 = in[1]? r1_2790 : r1_2789;
wire r2_1396;
assign r2_1396 = in[1]? r1_2792 : r1_2791;
wire r2_1397;
assign r2_1397 = in[1]? r1_2794 : r1_2793;
wire r2_1398;
assign r2_1398 = in[1]? r1_2796 : r1_2795;
wire r2_1399;
assign r2_1399 = in[1]? r1_2798 : r1_2797;
wire r2_1400;
assign r2_1400 = in[1]? r1_2800 : r1_2799;
wire r2_1401;
assign r2_1401 = in[1]? r1_2802 : r1_2801;
wire r2_1402;
assign r2_1402 = in[1]? r1_2804 : r1_2803;
wire r2_1403;
assign r2_1403 = in[1]? r1_2806 : r1_2805;
wire r2_1404;
assign r2_1404 = in[1]? r1_2808 : r1_2807;
wire r2_1405;
assign r2_1405 = in[1]? r1_2810 : r1_2809;
wire r2_1406;
assign r2_1406 = in[1]? r1_2812 : r1_2811;
wire r2_1407;
assign r2_1407 = in[1]? r1_2814 : r1_2813;
wire r2_1408;
assign r2_1408 = in[1]? r1_2816 : r1_2815;
wire r2_1409;
assign r2_1409 = in[1]? r1_2818 : r1_2817;
wire r2_1410;
assign r2_1410 = in[1]? r1_2820 : r1_2819;
wire r2_1411;
assign r2_1411 = in[1]? r1_2822 : r1_2821;
wire r2_1412;
assign r2_1412 = in[1]? r1_2824 : r1_2823;
wire r2_1413;
assign r2_1413 = in[1]? r1_2826 : r1_2825;
wire r2_1414;
assign r2_1414 = in[1]? r1_2828 : r1_2827;
wire r2_1415;
assign r2_1415 = in[1]? r1_2830 : r1_2829;
wire r2_1416;
assign r2_1416 = in[1]? r1_2832 : r1_2831;
wire r2_1417;
assign r2_1417 = in[1]? r1_2834 : r1_2833;
wire r2_1418;
assign r2_1418 = in[1]? r1_2836 : r1_2835;
wire r2_1419;
assign r2_1419 = in[1]? r1_2838 : r1_2837;
wire r2_1420;
assign r2_1420 = in[1]? r1_2840 : r1_2839;
wire r2_1421;
assign r2_1421 = in[1]? r1_2842 : r1_2841;
wire r2_1422;
assign r2_1422 = in[1]? r1_2844 : r1_2843;
wire r2_1423;
assign r2_1423 = in[1]? r1_2846 : r1_2845;
wire r2_1424;
assign r2_1424 = in[1]? r1_2848 : r1_2847;
wire r2_1425;
assign r2_1425 = in[1]? r1_2850 : r1_2849;
wire r2_1426;
assign r2_1426 = in[1]? r1_2852 : r1_2851;
wire r2_1427;
assign r2_1427 = in[1]? r1_2854 : r1_2853;
wire r2_1428;
assign r2_1428 = in[1]? r1_2856 : r1_2855;
wire r2_1429;
assign r2_1429 = in[1]? r1_2858 : r1_2857;
wire r2_1430;
assign r2_1430 = in[1]? r1_2860 : r1_2859;
wire r2_1431;
assign r2_1431 = in[1]? r1_2862 : r1_2861;
wire r2_1432;
assign r2_1432 = in[1]? r1_2864 : r1_2863;
wire r2_1433;
assign r2_1433 = in[1]? r1_2866 : r1_2865;
wire r2_1434;
assign r2_1434 = in[1]? r1_2868 : r1_2867;
wire r2_1435;
assign r2_1435 = in[1]? r1_2870 : r1_2869;
wire r2_1436;
assign r2_1436 = in[1]? r1_2872 : r1_2871;
wire r2_1437;
assign r2_1437 = in[1]? r1_2874 : r1_2873;
wire r2_1438;
assign r2_1438 = in[1]? r1_2876 : r1_2875;
wire r2_1439;
assign r2_1439 = in[1]? r1_2878 : r1_2877;
wire r2_1440;
assign r2_1440 = in[1]? r1_2880 : r1_2879;
wire r2_1441;
assign r2_1441 = in[1]? r1_2882 : r1_2881;
wire r2_1442;
assign r2_1442 = in[1]? r1_2884 : r1_2883;
wire r2_1443;
assign r2_1443 = in[1]? r1_2886 : r1_2885;
wire r2_1444;
assign r2_1444 = in[1]? r1_2888 : r1_2887;
wire r2_1445;
assign r2_1445 = in[1]? r1_2890 : r1_2889;
wire r2_1446;
assign r2_1446 = in[1]? r1_2892 : r1_2891;
wire r2_1447;
assign r2_1447 = in[1]? r1_2894 : r1_2893;
wire r2_1448;
assign r2_1448 = in[1]? r1_2896 : r1_2895;
wire r2_1449;
assign r2_1449 = in[1]? r1_2898 : r1_2897;
wire r2_1450;
assign r2_1450 = in[1]? r1_2900 : r1_2899;
wire r2_1451;
assign r2_1451 = in[1]? r1_2902 : r1_2901;
wire r2_1452;
assign r2_1452 = in[1]? r1_2904 : r1_2903;
wire r2_1453;
assign r2_1453 = in[1]? r1_2906 : r1_2905;
wire r2_1454;
assign r2_1454 = in[1]? r1_2908 : r1_2907;
wire r2_1455;
assign r2_1455 = in[1]? r1_2910 : r1_2909;
wire r2_1456;
assign r2_1456 = in[1]? r1_2912 : r1_2911;
wire r2_1457;
assign r2_1457 = in[1]? r1_2914 : r1_2913;
wire r2_1458;
assign r2_1458 = in[1]? r1_2916 : r1_2915;
wire r2_1459;
assign r2_1459 = in[1]? r1_2918 : r1_2917;
wire r2_1460;
assign r2_1460 = in[1]? r1_2920 : r1_2919;
wire r2_1461;
assign r2_1461 = in[1]? r1_2922 : r1_2921;
wire r2_1462;
assign r2_1462 = in[1]? r1_2924 : r1_2923;
wire r2_1463;
assign r2_1463 = in[1]? r1_2926 : r1_2925;
wire r2_1464;
assign r2_1464 = in[1]? r1_2928 : r1_2927;
wire r2_1465;
assign r2_1465 = in[1]? r1_2930 : r1_2929;
wire r2_1466;
assign r2_1466 = in[1]? r1_2932 : r1_2931;
wire r2_1467;
assign r2_1467 = in[1]? r1_2934 : r1_2933;
wire r2_1468;
assign r2_1468 = in[1]? r1_2936 : r1_2935;
wire r2_1469;
assign r2_1469 = in[1]? r1_2938 : r1_2937;
wire r2_1470;
assign r2_1470 = in[1]? r1_2940 : r1_2939;
wire r2_1471;
assign r2_1471 = in[1]? r1_2942 : r1_2941;
wire r2_1472;
assign r2_1472 = in[1]? r1_2944 : r1_2943;
wire r2_1473;
assign r2_1473 = in[1]? r1_2946 : r1_2945;
wire r2_1474;
assign r2_1474 = in[1]? r1_2948 : r1_2947;
wire r2_1475;
assign r2_1475 = in[1]? r1_2950 : r1_2949;
wire r2_1476;
assign r2_1476 = in[1]? r1_2952 : r1_2951;
wire r2_1477;
assign r2_1477 = in[1]? r1_2954 : r1_2953;
wire r2_1478;
assign r2_1478 = in[1]? r1_2956 : r1_2955;
wire r2_1479;
assign r2_1479 = in[1]? r1_2958 : r1_2957;
wire r2_1480;
assign r2_1480 = in[1]? r1_2960 : r1_2959;
wire r2_1481;
assign r2_1481 = in[1]? r1_2962 : r1_2961;
wire r2_1482;
assign r2_1482 = in[1]? r1_2964 : r1_2963;
wire r2_1483;
assign r2_1483 = in[1]? r1_2966 : r1_2965;
wire r2_1484;
assign r2_1484 = in[1]? r1_2968 : r1_2967;
wire r2_1485;
assign r2_1485 = in[1]? r1_2970 : r1_2969;
wire r2_1486;
assign r2_1486 = in[1]? r1_2972 : r1_2971;
wire r2_1487;
assign r2_1487 = in[1]? r1_2974 : r1_2973;
wire r2_1488;
assign r2_1488 = in[1]? r1_2976 : r1_2975;
wire r2_1489;
assign r2_1489 = in[1]? r1_2978 : r1_2977;
wire r2_1490;
assign r2_1490 = in[1]? r1_2980 : r1_2979;
wire r2_1491;
assign r2_1491 = in[1]? r1_2982 : r1_2981;
wire r2_1492;
assign r2_1492 = in[1]? r1_2984 : r1_2983;
wire r2_1493;
assign r2_1493 = in[1]? r1_2986 : r1_2985;
wire r2_1494;
assign r2_1494 = in[1]? r1_2988 : r1_2987;
wire r2_1495;
assign r2_1495 = in[1]? r1_2990 : r1_2989;
wire r2_1496;
assign r2_1496 = in[1]? r1_2992 : r1_2991;
wire r2_1497;
assign r2_1497 = in[1]? r1_2994 : r1_2993;
wire r2_1498;
assign r2_1498 = in[1]? r1_2996 : r1_2995;
wire r2_1499;
assign r2_1499 = in[1]? r1_2998 : r1_2997;
wire r2_1500;
assign r2_1500 = in[1]? r1_3000 : r1_2999;
wire r2_1501;
assign r2_1501 = in[1]? r1_3002 : r1_3001;
wire r2_1502;
assign r2_1502 = in[1]? r1_3004 : r1_3003;
wire r2_1503;
assign r2_1503 = in[1]? r1_3006 : r1_3005;
wire r2_1504;
assign r2_1504 = in[1]? r1_3008 : r1_3007;
wire r2_1505;
assign r2_1505 = in[1]? r1_3010 : r1_3009;
wire r2_1506;
assign r2_1506 = in[1]? r1_3012 : r1_3011;
wire r2_1507;
assign r2_1507 = in[1]? r1_3014 : r1_3013;
wire r2_1508;
assign r2_1508 = in[1]? r1_3016 : r1_3015;
wire r2_1509;
assign r2_1509 = in[1]? r1_3018 : r1_3017;
wire r2_1510;
assign r2_1510 = in[1]? r1_3020 : r1_3019;
wire r2_1511;
assign r2_1511 = in[1]? r1_3022 : r1_3021;
wire r2_1512;
assign r2_1512 = in[1]? r1_3024 : r1_3023;
wire r2_1513;
assign r2_1513 = in[1]? r1_3026 : r1_3025;
wire r2_1514;
assign r2_1514 = in[1]? r1_3028 : r1_3027;
wire r2_1515;
assign r2_1515 = in[1]? r1_3030 : r1_3029;
wire r2_1516;
assign r2_1516 = in[1]? r1_3032 : r1_3031;
wire r2_1517;
assign r2_1517 = in[1]? r1_3034 : r1_3033;
wire r2_1518;
assign r2_1518 = in[1]? r1_3036 : r1_3035;
wire r2_1519;
assign r2_1519 = in[1]? r1_3038 : r1_3037;
wire r2_1520;
assign r2_1520 = in[1]? r1_3040 : r1_3039;
wire r2_1521;
assign r2_1521 = in[1]? r1_3042 : r1_3041;
wire r2_1522;
assign r2_1522 = in[1]? r1_3044 : r1_3043;
wire r2_1523;
assign r2_1523 = in[1]? r1_3046 : r1_3045;
wire r2_1524;
assign r2_1524 = in[1]? r1_3048 : r1_3047;
wire r2_1525;
assign r2_1525 = in[1]? r1_3050 : r1_3049;
wire r2_1526;
assign r2_1526 = in[1]? r1_3052 : r1_3051;
wire r2_1527;
assign r2_1527 = in[1]? r1_3054 : r1_3053;
wire r2_1528;
assign r2_1528 = in[1]? r1_3056 : r1_3055;
wire r2_1529;
assign r2_1529 = in[1]? r1_3058 : r1_3057;
wire r2_1530;
assign r2_1530 = in[1]? r1_3060 : r1_3059;
wire r2_1531;
assign r2_1531 = in[1]? r1_3062 : r1_3061;
wire r2_1532;
assign r2_1532 = in[1]? r1_3064 : r1_3063;
wire r2_1533;
assign r2_1533 = in[1]? r1_3066 : r1_3065;
wire r2_1534;
assign r2_1534 = in[1]? r1_3068 : r1_3067;
wire r2_1535;
assign r2_1535 = in[1]? r1_3070 : r1_3069;
wire r2_1536;
assign r2_1536 = in[1]? r1_3072 : r1_3071;
wire r3_1;
assign r3_1 = in[2]? r2_2 : r2_1;
wire r3_2;
assign r3_2 = in[2]? r2_4 : r2_3;
wire r3_3;
assign r3_3 = in[2]? r2_6 : r2_5;
wire r3_4;
assign r3_4 = in[2]? r2_8 : r2_7;
wire r3_5;
assign r3_5 = in[2]? r2_10 : r2_9;
wire r3_6;
assign r3_6 = in[2]? r2_12 : r2_11;
wire r3_7;
assign r3_7 = in[2]? r2_14 : r2_13;
wire r3_8;
assign r3_8 = in[2]? r2_16 : r2_15;
wire r3_9;
assign r3_9 = in[2]? r2_18 : r2_17;
wire r3_10;
assign r3_10 = in[2]? r2_20 : r2_19;
wire r3_11;
assign r3_11 = in[2]? r2_22 : r2_21;
wire r3_12;
assign r3_12 = in[2]? r2_24 : r2_23;
wire r3_13;
assign r3_13 = in[2]? r2_26 : r2_25;
wire r3_14;
assign r3_14 = in[2]? r2_28 : r2_27;
wire r3_15;
assign r3_15 = in[2]? r2_30 : r2_29;
wire r3_16;
assign r3_16 = in[2]? r2_32 : r2_31;
wire r3_17;
assign r3_17 = in[2]? r2_34 : r2_33;
wire r3_18;
assign r3_18 = in[2]? r2_36 : r2_35;
wire r3_19;
assign r3_19 = in[2]? r2_38 : r2_37;
wire r3_20;
assign r3_20 = in[2]? r2_40 : r2_39;
wire r3_21;
assign r3_21 = in[2]? r2_42 : r2_41;
wire r3_22;
assign r3_22 = in[2]? r2_44 : r2_43;
wire r3_23;
assign r3_23 = in[2]? r2_46 : r2_45;
wire r3_24;
assign r3_24 = in[2]? r2_48 : r2_47;
wire r3_25;
assign r3_25 = in[2]? r2_50 : r2_49;
wire r3_26;
assign r3_26 = in[2]? r2_52 : r2_51;
wire r3_27;
assign r3_27 = in[2]? r2_54 : r2_53;
wire r3_28;
assign r3_28 = in[2]? r2_56 : r2_55;
wire r3_29;
assign r3_29 = in[2]? r2_58 : r2_57;
wire r3_30;
assign r3_30 = in[2]? r2_60 : r2_59;
wire r3_31;
assign r3_31 = in[2]? r2_62 : r2_61;
wire r3_32;
assign r3_32 = in[2]? r2_64 : r2_63;
wire r3_33;
assign r3_33 = in[2]? r2_66 : r2_65;
wire r3_34;
assign r3_34 = in[2]? r2_68 : r2_67;
wire r3_35;
assign r3_35 = in[2]? r2_70 : r2_69;
wire r3_36;
assign r3_36 = in[2]? r2_72 : r2_71;
wire r3_37;
assign r3_37 = in[2]? r2_74 : r2_73;
wire r3_38;
assign r3_38 = in[2]? r2_76 : r2_75;
wire r3_39;
assign r3_39 = in[2]? r2_78 : r2_77;
wire r3_40;
assign r3_40 = in[2]? r2_80 : r2_79;
wire r3_41;
assign r3_41 = in[2]? r2_82 : r2_81;
wire r3_42;
assign r3_42 = in[2]? r2_84 : r2_83;
wire r3_43;
assign r3_43 = in[2]? r2_86 : r2_85;
wire r3_44;
assign r3_44 = in[2]? r2_88 : r2_87;
wire r3_45;
assign r3_45 = in[2]? r2_90 : r2_89;
wire r3_46;
assign r3_46 = in[2]? r2_92 : r2_91;
wire r3_47;
assign r3_47 = in[2]? r2_94 : r2_93;
wire r3_48;
assign r3_48 = in[2]? r2_96 : r2_95;
wire r3_49;
assign r3_49 = in[2]? r2_98 : r2_97;
wire r3_50;
assign r3_50 = in[2]? r2_100 : r2_99;
wire r3_51;
assign r3_51 = in[2]? r2_102 : r2_101;
wire r3_52;
assign r3_52 = in[2]? r2_104 : r2_103;
wire r3_53;
assign r3_53 = in[2]? r2_106 : r2_105;
wire r3_54;
assign r3_54 = in[2]? r2_108 : r2_107;
wire r3_55;
assign r3_55 = in[2]? r2_110 : r2_109;
wire r3_56;
assign r3_56 = in[2]? r2_112 : r2_111;
wire r3_57;
assign r3_57 = in[2]? r2_114 : r2_113;
wire r3_58;
assign r3_58 = in[2]? r2_116 : r2_115;
wire r3_59;
assign r3_59 = in[2]? r2_118 : r2_117;
wire r3_60;
assign r3_60 = in[2]? r2_120 : r2_119;
wire r3_61;
assign r3_61 = in[2]? r2_122 : r2_121;
wire r3_62;
assign r3_62 = in[2]? r2_124 : r2_123;
wire r3_63;
assign r3_63 = in[2]? r2_126 : r2_125;
wire r3_64;
assign r3_64 = in[2]? r2_128 : r2_127;
wire r3_65;
assign r3_65 = in[2]? r2_130 : r2_129;
wire r3_66;
assign r3_66 = in[2]? r2_132 : r2_131;
wire r3_67;
assign r3_67 = in[2]? r2_134 : r2_133;
wire r3_68;
assign r3_68 = in[2]? r2_136 : r2_135;
wire r3_69;
assign r3_69 = in[2]? r2_138 : r2_137;
wire r3_70;
assign r3_70 = in[2]? r2_140 : r2_139;
wire r3_71;
assign r3_71 = in[2]? r2_142 : r2_141;
wire r3_72;
assign r3_72 = in[2]? r2_144 : r2_143;
wire r3_73;
assign r3_73 = in[2]? r2_146 : r2_145;
wire r3_74;
assign r3_74 = in[2]? r2_148 : r2_147;
wire r3_75;
assign r3_75 = in[2]? r2_150 : r2_149;
wire r3_76;
assign r3_76 = in[2]? r2_152 : r2_151;
wire r3_77;
assign r3_77 = in[2]? r2_154 : r2_153;
wire r3_78;
assign r3_78 = in[2]? r2_156 : r2_155;
wire r3_79;
assign r3_79 = in[2]? r2_158 : r2_157;
wire r3_80;
assign r3_80 = in[2]? r2_160 : r2_159;
wire r3_81;
assign r3_81 = in[2]? r2_162 : r2_161;
wire r3_82;
assign r3_82 = in[2]? r2_164 : r2_163;
wire r3_83;
assign r3_83 = in[2]? r2_166 : r2_165;
wire r3_84;
assign r3_84 = in[2]? r2_168 : r2_167;
wire r3_85;
assign r3_85 = in[2]? r2_170 : r2_169;
wire r3_86;
assign r3_86 = in[2]? r2_172 : r2_171;
wire r3_87;
assign r3_87 = in[2]? r2_174 : r2_173;
wire r3_88;
assign r3_88 = in[2]? r2_176 : r2_175;
wire r3_89;
assign r3_89 = in[2]? r2_178 : r2_177;
wire r3_90;
assign r3_90 = in[2]? r2_180 : r2_179;
wire r3_91;
assign r3_91 = in[2]? r2_182 : r2_181;
wire r3_92;
assign r3_92 = in[2]? r2_184 : r2_183;
wire r3_93;
assign r3_93 = in[2]? r2_186 : r2_185;
wire r3_94;
assign r3_94 = in[2]? r2_188 : r2_187;
wire r3_95;
assign r3_95 = in[2]? r2_190 : r2_189;
wire r3_96;
assign r3_96 = in[2]? r2_192 : r2_191;
wire r3_97;
assign r3_97 = in[2]? r2_194 : r2_193;
wire r3_98;
assign r3_98 = in[2]? r2_196 : r2_195;
wire r3_99;
assign r3_99 = in[2]? r2_198 : r2_197;
wire r3_100;
assign r3_100 = in[2]? r2_200 : r2_199;
wire r3_101;
assign r3_101 = in[2]? r2_202 : r2_201;
wire r3_102;
assign r3_102 = in[2]? r2_204 : r2_203;
wire r3_103;
assign r3_103 = in[2]? r2_206 : r2_205;
wire r3_104;
assign r3_104 = in[2]? r2_208 : r2_207;
wire r3_105;
assign r3_105 = in[2]? r2_210 : r2_209;
wire r3_106;
assign r3_106 = in[2]? r2_212 : r2_211;
wire r3_107;
assign r3_107 = in[2]? r2_214 : r2_213;
wire r3_108;
assign r3_108 = in[2]? r2_216 : r2_215;
wire r3_109;
assign r3_109 = in[2]? r2_218 : r2_217;
wire r3_110;
assign r3_110 = in[2]? r2_220 : r2_219;
wire r3_111;
assign r3_111 = in[2]? r2_222 : r2_221;
wire r3_112;
assign r3_112 = in[2]? r2_224 : r2_223;
wire r3_113;
assign r3_113 = in[2]? r2_226 : r2_225;
wire r3_114;
assign r3_114 = in[2]? r2_228 : r2_227;
wire r3_115;
assign r3_115 = in[2]? r2_230 : r2_229;
wire r3_116;
assign r3_116 = in[2]? r2_232 : r2_231;
wire r3_117;
assign r3_117 = in[2]? r2_234 : r2_233;
wire r3_118;
assign r3_118 = in[2]? r2_236 : r2_235;
wire r3_119;
assign r3_119 = in[2]? r2_238 : r2_237;
wire r3_120;
assign r3_120 = in[2]? r2_240 : r2_239;
wire r3_121;
assign r3_121 = in[2]? r2_242 : r2_241;
wire r3_122;
assign r3_122 = in[2]? r2_244 : r2_243;
wire r3_123;
assign r3_123 = in[2]? r2_246 : r2_245;
wire r3_124;
assign r3_124 = in[2]? r2_248 : r2_247;
wire r3_125;
assign r3_125 = in[2]? r2_250 : r2_249;
wire r3_126;
assign r3_126 = in[2]? r2_252 : r2_251;
wire r3_127;
assign r3_127 = in[2]? r2_254 : r2_253;
wire r3_128;
assign r3_128 = in[2]? r2_256 : r2_255;
wire r3_129;
assign r3_129 = in[2]? r2_258 : r2_257;
wire r3_130;
assign r3_130 = in[2]? r2_260 : r2_259;
wire r3_131;
assign r3_131 = in[2]? r2_262 : r2_261;
wire r3_132;
assign r3_132 = in[2]? r2_264 : r2_263;
wire r3_133;
assign r3_133 = in[2]? r2_266 : r2_265;
wire r3_134;
assign r3_134 = in[2]? r2_268 : r2_267;
wire r3_135;
assign r3_135 = in[2]? r2_270 : r2_269;
wire r3_136;
assign r3_136 = in[2]? r2_272 : r2_271;
wire r3_137;
assign r3_137 = in[2]? r2_274 : r2_273;
wire r3_138;
assign r3_138 = in[2]? r2_276 : r2_275;
wire r3_139;
assign r3_139 = in[2]? r2_278 : r2_277;
wire r3_140;
assign r3_140 = in[2]? r2_280 : r2_279;
wire r3_141;
assign r3_141 = in[2]? r2_282 : r2_281;
wire r3_142;
assign r3_142 = in[2]? r2_284 : r2_283;
wire r3_143;
assign r3_143 = in[2]? r2_286 : r2_285;
wire r3_144;
assign r3_144 = in[2]? r2_288 : r2_287;
wire r3_145;
assign r3_145 = in[2]? r2_290 : r2_289;
wire r3_146;
assign r3_146 = in[2]? r2_292 : r2_291;
wire r3_147;
assign r3_147 = in[2]? r2_294 : r2_293;
wire r3_148;
assign r3_148 = in[2]? r2_296 : r2_295;
wire r3_149;
assign r3_149 = in[2]? r2_298 : r2_297;
wire r3_150;
assign r3_150 = in[2]? r2_300 : r2_299;
wire r3_151;
assign r3_151 = in[2]? r2_302 : r2_301;
wire r3_152;
assign r3_152 = in[2]? r2_304 : r2_303;
wire r3_153;
assign r3_153 = in[2]? r2_306 : r2_305;
wire r3_154;
assign r3_154 = in[2]? r2_308 : r2_307;
wire r3_155;
assign r3_155 = in[2]? r2_310 : r2_309;
wire r3_156;
assign r3_156 = in[2]? r2_312 : r2_311;
wire r3_157;
assign r3_157 = in[2]? r2_314 : r2_313;
wire r3_158;
assign r3_158 = in[2]? r2_316 : r2_315;
wire r3_159;
assign r3_159 = in[2]? r2_318 : r2_317;
wire r3_160;
assign r3_160 = in[2]? r2_320 : r2_319;
wire r3_161;
assign r3_161 = in[2]? r2_322 : r2_321;
wire r3_162;
assign r3_162 = in[2]? r2_324 : r2_323;
wire r3_163;
assign r3_163 = in[2]? r2_326 : r2_325;
wire r3_164;
assign r3_164 = in[2]? r2_328 : r2_327;
wire r3_165;
assign r3_165 = in[2]? r2_330 : r2_329;
wire r3_166;
assign r3_166 = in[2]? r2_332 : r2_331;
wire r3_167;
assign r3_167 = in[2]? r2_334 : r2_333;
wire r3_168;
assign r3_168 = in[2]? r2_336 : r2_335;
wire r3_169;
assign r3_169 = in[2]? r2_338 : r2_337;
wire r3_170;
assign r3_170 = in[2]? r2_340 : r2_339;
wire r3_171;
assign r3_171 = in[2]? r2_342 : r2_341;
wire r3_172;
assign r3_172 = in[2]? r2_344 : r2_343;
wire r3_173;
assign r3_173 = in[2]? r2_346 : r2_345;
wire r3_174;
assign r3_174 = in[2]? r2_348 : r2_347;
wire r3_175;
assign r3_175 = in[2]? r2_350 : r2_349;
wire r3_176;
assign r3_176 = in[2]? r2_352 : r2_351;
wire r3_177;
assign r3_177 = in[2]? r2_354 : r2_353;
wire r3_178;
assign r3_178 = in[2]? r2_356 : r2_355;
wire r3_179;
assign r3_179 = in[2]? r2_358 : r2_357;
wire r3_180;
assign r3_180 = in[2]? r2_360 : r2_359;
wire r3_181;
assign r3_181 = in[2]? r2_362 : r2_361;
wire r3_182;
assign r3_182 = in[2]? r2_364 : r2_363;
wire r3_183;
assign r3_183 = in[2]? r2_366 : r2_365;
wire r3_184;
assign r3_184 = in[2]? r2_368 : r2_367;
wire r3_185;
assign r3_185 = in[2]? r2_370 : r2_369;
wire r3_186;
assign r3_186 = in[2]? r2_372 : r2_371;
wire r3_187;
assign r3_187 = in[2]? r2_374 : r2_373;
wire r3_188;
assign r3_188 = in[2]? r2_376 : r2_375;
wire r3_189;
assign r3_189 = in[2]? r2_378 : r2_377;
wire r3_190;
assign r3_190 = in[2]? r2_380 : r2_379;
wire r3_191;
assign r3_191 = in[2]? r2_382 : r2_381;
wire r3_192;
assign r3_192 = in[2]? r2_384 : r2_383;
wire r3_193;
assign r3_193 = in[2]? r2_386 : r2_385;
wire r3_194;
assign r3_194 = in[2]? r2_388 : r2_387;
wire r3_195;
assign r3_195 = in[2]? r2_390 : r2_389;
wire r3_196;
assign r3_196 = in[2]? r2_392 : r2_391;
wire r3_197;
assign r3_197 = in[2]? r2_394 : r2_393;
wire r3_198;
assign r3_198 = in[2]? r2_396 : r2_395;
wire r3_199;
assign r3_199 = in[2]? r2_398 : r2_397;
wire r3_200;
assign r3_200 = in[2]? r2_400 : r2_399;
wire r3_201;
assign r3_201 = in[2]? r2_402 : r2_401;
wire r3_202;
assign r3_202 = in[2]? r2_404 : r2_403;
wire r3_203;
assign r3_203 = in[2]? r2_406 : r2_405;
wire r3_204;
assign r3_204 = in[2]? r2_408 : r2_407;
wire r3_205;
assign r3_205 = in[2]? r2_410 : r2_409;
wire r3_206;
assign r3_206 = in[2]? r2_412 : r2_411;
wire r3_207;
assign r3_207 = in[2]? r2_414 : r2_413;
wire r3_208;
assign r3_208 = in[2]? r2_416 : r2_415;
wire r3_209;
assign r3_209 = in[2]? r2_418 : r2_417;
wire r3_210;
assign r3_210 = in[2]? r2_420 : r2_419;
wire r3_211;
assign r3_211 = in[2]? r2_422 : r2_421;
wire r3_212;
assign r3_212 = in[2]? r2_424 : r2_423;
wire r3_213;
assign r3_213 = in[2]? r2_426 : r2_425;
wire r3_214;
assign r3_214 = in[2]? r2_428 : r2_427;
wire r3_215;
assign r3_215 = in[2]? r2_430 : r2_429;
wire r3_216;
assign r3_216 = in[2]? r2_432 : r2_431;
wire r3_217;
assign r3_217 = in[2]? r2_434 : r2_433;
wire r3_218;
assign r3_218 = in[2]? r2_436 : r2_435;
wire r3_219;
assign r3_219 = in[2]? r2_438 : r2_437;
wire r3_220;
assign r3_220 = in[2]? r2_440 : r2_439;
wire r3_221;
assign r3_221 = in[2]? r2_442 : r2_441;
wire r3_222;
assign r3_222 = in[2]? r2_444 : r2_443;
wire r3_223;
assign r3_223 = in[2]? r2_446 : r2_445;
wire r3_224;
assign r3_224 = in[2]? r2_448 : r2_447;
wire r3_225;
assign r3_225 = in[2]? r2_450 : r2_449;
wire r3_226;
assign r3_226 = in[2]? r2_452 : r2_451;
wire r3_227;
assign r3_227 = in[2]? r2_454 : r2_453;
wire r3_228;
assign r3_228 = in[2]? r2_456 : r2_455;
wire r3_229;
assign r3_229 = in[2]? r2_458 : r2_457;
wire r3_230;
assign r3_230 = in[2]? r2_460 : r2_459;
wire r3_231;
assign r3_231 = in[2]? r2_462 : r2_461;
wire r3_232;
assign r3_232 = in[2]? r2_464 : r2_463;
wire r3_233;
assign r3_233 = in[2]? r2_466 : r2_465;
wire r3_234;
assign r3_234 = in[2]? r2_468 : r2_467;
wire r3_235;
assign r3_235 = in[2]? r2_470 : r2_469;
wire r3_236;
assign r3_236 = in[2]? r2_472 : r2_471;
wire r3_237;
assign r3_237 = in[2]? r2_474 : r2_473;
wire r3_238;
assign r3_238 = in[2]? r2_476 : r2_475;
wire r3_239;
assign r3_239 = in[2]? r2_478 : r2_477;
wire r3_240;
assign r3_240 = in[2]? r2_480 : r2_479;
wire r3_241;
assign r3_241 = in[2]? r2_482 : r2_481;
wire r3_242;
assign r3_242 = in[2]? r2_484 : r2_483;
wire r3_243;
assign r3_243 = in[2]? r2_486 : r2_485;
wire r3_244;
assign r3_244 = in[2]? r2_488 : r2_487;
wire r3_245;
assign r3_245 = in[2]? r2_490 : r2_489;
wire r3_246;
assign r3_246 = in[2]? r2_492 : r2_491;
wire r3_247;
assign r3_247 = in[2]? r2_494 : r2_493;
wire r3_248;
assign r3_248 = in[2]? r2_496 : r2_495;
wire r3_249;
assign r3_249 = in[2]? r2_498 : r2_497;
wire r3_250;
assign r3_250 = in[2]? r2_500 : r2_499;
wire r3_251;
assign r3_251 = in[2]? r2_502 : r2_501;
wire r3_252;
assign r3_252 = in[2]? r2_504 : r2_503;
wire r3_253;
assign r3_253 = in[2]? r2_506 : r2_505;
wire r3_254;
assign r3_254 = in[2]? r2_508 : r2_507;
wire r3_255;
assign r3_255 = in[2]? r2_510 : r2_509;
wire r3_256;
assign r3_256 = in[2]? r2_512 : r2_511;
wire r3_257;
assign r3_257 = in[2]? r2_514 : r2_513;
wire r3_258;
assign r3_258 = in[2]? r2_516 : r2_515;
wire r3_259;
assign r3_259 = in[2]? r2_518 : r2_517;
wire r3_260;
assign r3_260 = in[2]? r2_520 : r2_519;
wire r3_261;
assign r3_261 = in[2]? r2_522 : r2_521;
wire r3_262;
assign r3_262 = in[2]? r2_524 : r2_523;
wire r3_263;
assign r3_263 = in[2]? r2_526 : r2_525;
wire r3_264;
assign r3_264 = in[2]? r2_528 : r2_527;
wire r3_265;
assign r3_265 = in[2]? r2_530 : r2_529;
wire r3_266;
assign r3_266 = in[2]? r2_532 : r2_531;
wire r3_267;
assign r3_267 = in[2]? r2_534 : r2_533;
wire r3_268;
assign r3_268 = in[2]? r2_536 : r2_535;
wire r3_269;
assign r3_269 = in[2]? r2_538 : r2_537;
wire r3_270;
assign r3_270 = in[2]? r2_540 : r2_539;
wire r3_271;
assign r3_271 = in[2]? r2_542 : r2_541;
wire r3_272;
assign r3_272 = in[2]? r2_544 : r2_543;
wire r3_273;
assign r3_273 = in[2]? r2_546 : r2_545;
wire r3_274;
assign r3_274 = in[2]? r2_548 : r2_547;
wire r3_275;
assign r3_275 = in[2]? r2_550 : r2_549;
wire r3_276;
assign r3_276 = in[2]? r2_552 : r2_551;
wire r3_277;
assign r3_277 = in[2]? r2_554 : r2_553;
wire r3_278;
assign r3_278 = in[2]? r2_556 : r2_555;
wire r3_279;
assign r3_279 = in[2]? r2_558 : r2_557;
wire r3_280;
assign r3_280 = in[2]? r2_560 : r2_559;
wire r3_281;
assign r3_281 = in[2]? r2_562 : r2_561;
wire r3_282;
assign r3_282 = in[2]? r2_564 : r2_563;
wire r3_283;
assign r3_283 = in[2]? r2_566 : r2_565;
wire r3_284;
assign r3_284 = in[2]? r2_568 : r2_567;
wire r3_285;
assign r3_285 = in[2]? r2_570 : r2_569;
wire r3_286;
assign r3_286 = in[2]? r2_572 : r2_571;
wire r3_287;
assign r3_287 = in[2]? r2_574 : r2_573;
wire r3_288;
assign r3_288 = in[2]? r2_576 : r2_575;
wire r3_289;
assign r3_289 = in[2]? r2_578 : r2_577;
wire r3_290;
assign r3_290 = in[2]? r2_580 : r2_579;
wire r3_291;
assign r3_291 = in[2]? r2_582 : r2_581;
wire r3_292;
assign r3_292 = in[2]? r2_584 : r2_583;
wire r3_293;
assign r3_293 = in[2]? r2_586 : r2_585;
wire r3_294;
assign r3_294 = in[2]? r2_588 : r2_587;
wire r3_295;
assign r3_295 = in[2]? r2_590 : r2_589;
wire r3_296;
assign r3_296 = in[2]? r2_592 : r2_591;
wire r3_297;
assign r3_297 = in[2]? r2_594 : r2_593;
wire r3_298;
assign r3_298 = in[2]? r2_596 : r2_595;
wire r3_299;
assign r3_299 = in[2]? r2_598 : r2_597;
wire r3_300;
assign r3_300 = in[2]? r2_600 : r2_599;
wire r3_301;
assign r3_301 = in[2]? r2_602 : r2_601;
wire r3_302;
assign r3_302 = in[2]? r2_604 : r2_603;
wire r3_303;
assign r3_303 = in[2]? r2_606 : r2_605;
wire r3_304;
assign r3_304 = in[2]? r2_608 : r2_607;
wire r3_305;
assign r3_305 = in[2]? r2_610 : r2_609;
wire r3_306;
assign r3_306 = in[2]? r2_612 : r2_611;
wire r3_307;
assign r3_307 = in[2]? r2_614 : r2_613;
wire r3_308;
assign r3_308 = in[2]? r2_616 : r2_615;
wire r3_309;
assign r3_309 = in[2]? r2_618 : r2_617;
wire r3_310;
assign r3_310 = in[2]? r2_620 : r2_619;
wire r3_311;
assign r3_311 = in[2]? r2_622 : r2_621;
wire r3_312;
assign r3_312 = in[2]? r2_624 : r2_623;
wire r3_313;
assign r3_313 = in[2]? r2_626 : r2_625;
wire r3_314;
assign r3_314 = in[2]? r2_628 : r2_627;
wire r3_315;
assign r3_315 = in[2]? r2_630 : r2_629;
wire r3_316;
assign r3_316 = in[2]? r2_632 : r2_631;
wire r3_317;
assign r3_317 = in[2]? r2_634 : r2_633;
wire r3_318;
assign r3_318 = in[2]? r2_636 : r2_635;
wire r3_319;
assign r3_319 = in[2]? r2_638 : r2_637;
wire r3_320;
assign r3_320 = in[2]? r2_640 : r2_639;
wire r3_321;
assign r3_321 = in[2]? r2_642 : r2_641;
wire r3_322;
assign r3_322 = in[2]? r2_644 : r2_643;
wire r3_323;
assign r3_323 = in[2]? r2_646 : r2_645;
wire r3_324;
assign r3_324 = in[2]? r2_648 : r2_647;
wire r3_325;
assign r3_325 = in[2]? r2_650 : r2_649;
wire r3_326;
assign r3_326 = in[2]? r2_652 : r2_651;
wire r3_327;
assign r3_327 = in[2]? r2_654 : r2_653;
wire r3_328;
assign r3_328 = in[2]? r2_656 : r2_655;
wire r3_329;
assign r3_329 = in[2]? r2_658 : r2_657;
wire r3_330;
assign r3_330 = in[2]? r2_660 : r2_659;
wire r3_331;
assign r3_331 = in[2]? r2_662 : r2_661;
wire r3_332;
assign r3_332 = in[2]? r2_664 : r2_663;
wire r3_333;
assign r3_333 = in[2]? r2_666 : r2_665;
wire r3_334;
assign r3_334 = in[2]? r2_668 : r2_667;
wire r3_335;
assign r3_335 = in[2]? r2_670 : r2_669;
wire r3_336;
assign r3_336 = in[2]? r2_672 : r2_671;
wire r3_337;
assign r3_337 = in[2]? r2_674 : r2_673;
wire r3_338;
assign r3_338 = in[2]? r2_676 : r2_675;
wire r3_339;
assign r3_339 = in[2]? r2_678 : r2_677;
wire r3_340;
assign r3_340 = in[2]? r2_680 : r2_679;
wire r3_341;
assign r3_341 = in[2]? r2_682 : r2_681;
wire r3_342;
assign r3_342 = in[2]? r2_684 : r2_683;
wire r3_343;
assign r3_343 = in[2]? r2_686 : r2_685;
wire r3_344;
assign r3_344 = in[2]? r2_688 : r2_687;
wire r3_345;
assign r3_345 = in[2]? r2_690 : r2_689;
wire r3_346;
assign r3_346 = in[2]? r2_692 : r2_691;
wire r3_347;
assign r3_347 = in[2]? r2_694 : r2_693;
wire r3_348;
assign r3_348 = in[2]? r2_696 : r2_695;
wire r3_349;
assign r3_349 = in[2]? r2_698 : r2_697;
wire r3_350;
assign r3_350 = in[2]? r2_700 : r2_699;
wire r3_351;
assign r3_351 = in[2]? r2_702 : r2_701;
wire r3_352;
assign r3_352 = in[2]? r2_704 : r2_703;
wire r3_353;
assign r3_353 = in[2]? r2_706 : r2_705;
wire r3_354;
assign r3_354 = in[2]? r2_708 : r2_707;
wire r3_355;
assign r3_355 = in[2]? r2_710 : r2_709;
wire r3_356;
assign r3_356 = in[2]? r2_712 : r2_711;
wire r3_357;
assign r3_357 = in[2]? r2_714 : r2_713;
wire r3_358;
assign r3_358 = in[2]? r2_716 : r2_715;
wire r3_359;
assign r3_359 = in[2]? r2_718 : r2_717;
wire r3_360;
assign r3_360 = in[2]? r2_720 : r2_719;
wire r3_361;
assign r3_361 = in[2]? r2_722 : r2_721;
wire r3_362;
assign r3_362 = in[2]? r2_724 : r2_723;
wire r3_363;
assign r3_363 = in[2]? r2_726 : r2_725;
wire r3_364;
assign r3_364 = in[2]? r2_728 : r2_727;
wire r3_365;
assign r3_365 = in[2]? r2_730 : r2_729;
wire r3_366;
assign r3_366 = in[2]? r2_732 : r2_731;
wire r3_367;
assign r3_367 = in[2]? r2_734 : r2_733;
wire r3_368;
assign r3_368 = in[2]? r2_736 : r2_735;
wire r3_369;
assign r3_369 = in[2]? r2_738 : r2_737;
wire r3_370;
assign r3_370 = in[2]? r2_740 : r2_739;
wire r3_371;
assign r3_371 = in[2]? r2_742 : r2_741;
wire r3_372;
assign r3_372 = in[2]? r2_744 : r2_743;
wire r3_373;
assign r3_373 = in[2]? r2_746 : r2_745;
wire r3_374;
assign r3_374 = in[2]? r2_748 : r2_747;
wire r3_375;
assign r3_375 = in[2]? r2_750 : r2_749;
wire r3_376;
assign r3_376 = in[2]? r2_752 : r2_751;
wire r3_377;
assign r3_377 = in[2]? r2_754 : r2_753;
wire r3_378;
assign r3_378 = in[2]? r2_756 : r2_755;
wire r3_379;
assign r3_379 = in[2]? r2_758 : r2_757;
wire r3_380;
assign r3_380 = in[2]? r2_760 : r2_759;
wire r3_381;
assign r3_381 = in[2]? r2_762 : r2_761;
wire r3_382;
assign r3_382 = in[2]? r2_764 : r2_763;
wire r3_383;
assign r3_383 = in[2]? r2_766 : r2_765;
wire r3_384;
assign r3_384 = in[2]? r2_768 : r2_767;
wire r3_385;
assign r3_385 = in[2]? r2_770 : r2_769;
wire r3_386;
assign r3_386 = in[2]? r2_772 : r2_771;
wire r3_387;
assign r3_387 = in[2]? r2_774 : r2_773;
wire r3_388;
assign r3_388 = in[2]? r2_776 : r2_775;
wire r3_389;
assign r3_389 = in[2]? r2_778 : r2_777;
wire r3_390;
assign r3_390 = in[2]? r2_780 : r2_779;
wire r3_391;
assign r3_391 = in[2]? r2_782 : r2_781;
wire r3_392;
assign r3_392 = in[2]? r2_784 : r2_783;
wire r3_393;
assign r3_393 = in[2]? r2_786 : r2_785;
wire r3_394;
assign r3_394 = in[2]? r2_788 : r2_787;
wire r3_395;
assign r3_395 = in[2]? r2_790 : r2_789;
wire r3_396;
assign r3_396 = in[2]? r2_792 : r2_791;
wire r3_397;
assign r3_397 = in[2]? r2_794 : r2_793;
wire r3_398;
assign r3_398 = in[2]? r2_796 : r2_795;
wire r3_399;
assign r3_399 = in[2]? r2_798 : r2_797;
wire r3_400;
assign r3_400 = in[2]? r2_800 : r2_799;
wire r3_401;
assign r3_401 = in[2]? r2_802 : r2_801;
wire r3_402;
assign r3_402 = in[2]? r2_804 : r2_803;
wire r3_403;
assign r3_403 = in[2]? r2_806 : r2_805;
wire r3_404;
assign r3_404 = in[2]? r2_808 : r2_807;
wire r3_405;
assign r3_405 = in[2]? r2_810 : r2_809;
wire r3_406;
assign r3_406 = in[2]? r2_812 : r2_811;
wire r3_407;
assign r3_407 = in[2]? r2_814 : r2_813;
wire r3_408;
assign r3_408 = in[2]? r2_816 : r2_815;
wire r3_409;
assign r3_409 = in[2]? r2_818 : r2_817;
wire r3_410;
assign r3_410 = in[2]? r2_820 : r2_819;
wire r3_411;
assign r3_411 = in[2]? r2_822 : r2_821;
wire r3_412;
assign r3_412 = in[2]? r2_824 : r2_823;
wire r3_413;
assign r3_413 = in[2]? r2_826 : r2_825;
wire r3_414;
assign r3_414 = in[2]? r2_828 : r2_827;
wire r3_415;
assign r3_415 = in[2]? r2_830 : r2_829;
wire r3_416;
assign r3_416 = in[2]? r2_832 : r2_831;
wire r3_417;
assign r3_417 = in[2]? r2_834 : r2_833;
wire r3_418;
assign r3_418 = in[2]? r2_836 : r2_835;
wire r3_419;
assign r3_419 = in[2]? r2_838 : r2_837;
wire r3_420;
assign r3_420 = in[2]? r2_840 : r2_839;
wire r3_421;
assign r3_421 = in[2]? r2_842 : r2_841;
wire r3_422;
assign r3_422 = in[2]? r2_844 : r2_843;
wire r3_423;
assign r3_423 = in[2]? r2_846 : r2_845;
wire r3_424;
assign r3_424 = in[2]? r2_848 : r2_847;
wire r3_425;
assign r3_425 = in[2]? r2_850 : r2_849;
wire r3_426;
assign r3_426 = in[2]? r2_852 : r2_851;
wire r3_427;
assign r3_427 = in[2]? r2_854 : r2_853;
wire r3_428;
assign r3_428 = in[2]? r2_856 : r2_855;
wire r3_429;
assign r3_429 = in[2]? r2_858 : r2_857;
wire r3_430;
assign r3_430 = in[2]? r2_860 : r2_859;
wire r3_431;
assign r3_431 = in[2]? r2_862 : r2_861;
wire r3_432;
assign r3_432 = in[2]? r2_864 : r2_863;
wire r3_433;
assign r3_433 = in[2]? r2_866 : r2_865;
wire r3_434;
assign r3_434 = in[2]? r2_868 : r2_867;
wire r3_435;
assign r3_435 = in[2]? r2_870 : r2_869;
wire r3_436;
assign r3_436 = in[2]? r2_872 : r2_871;
wire r3_437;
assign r3_437 = in[2]? r2_874 : r2_873;
wire r3_438;
assign r3_438 = in[2]? r2_876 : r2_875;
wire r3_439;
assign r3_439 = in[2]? r2_878 : r2_877;
wire r3_440;
assign r3_440 = in[2]? r2_880 : r2_879;
wire r3_441;
assign r3_441 = in[2]? r2_882 : r2_881;
wire r3_442;
assign r3_442 = in[2]? r2_884 : r2_883;
wire r3_443;
assign r3_443 = in[2]? r2_886 : r2_885;
wire r3_444;
assign r3_444 = in[2]? r2_888 : r2_887;
wire r3_445;
assign r3_445 = in[2]? r2_890 : r2_889;
wire r3_446;
assign r3_446 = in[2]? r2_892 : r2_891;
wire r3_447;
assign r3_447 = in[2]? r2_894 : r2_893;
wire r3_448;
assign r3_448 = in[2]? r2_896 : r2_895;
wire r3_449;
assign r3_449 = in[2]? r2_898 : r2_897;
wire r3_450;
assign r3_450 = in[2]? r2_900 : r2_899;
wire r3_451;
assign r3_451 = in[2]? r2_902 : r2_901;
wire r3_452;
assign r3_452 = in[2]? r2_904 : r2_903;
wire r3_453;
assign r3_453 = in[2]? r2_906 : r2_905;
wire r3_454;
assign r3_454 = in[2]? r2_908 : r2_907;
wire r3_455;
assign r3_455 = in[2]? r2_910 : r2_909;
wire r3_456;
assign r3_456 = in[2]? r2_912 : r2_911;
wire r3_457;
assign r3_457 = in[2]? r2_914 : r2_913;
wire r3_458;
assign r3_458 = in[2]? r2_916 : r2_915;
wire r3_459;
assign r3_459 = in[2]? r2_918 : r2_917;
wire r3_460;
assign r3_460 = in[2]? r2_920 : r2_919;
wire r3_461;
assign r3_461 = in[2]? r2_922 : r2_921;
wire r3_462;
assign r3_462 = in[2]? r2_924 : r2_923;
wire r3_463;
assign r3_463 = in[2]? r2_926 : r2_925;
wire r3_464;
assign r3_464 = in[2]? r2_928 : r2_927;
wire r3_465;
assign r3_465 = in[2]? r2_930 : r2_929;
wire r3_466;
assign r3_466 = in[2]? r2_932 : r2_931;
wire r3_467;
assign r3_467 = in[2]? r2_934 : r2_933;
wire r3_468;
assign r3_468 = in[2]? r2_936 : r2_935;
wire r3_469;
assign r3_469 = in[2]? r2_938 : r2_937;
wire r3_470;
assign r3_470 = in[2]? r2_940 : r2_939;
wire r3_471;
assign r3_471 = in[2]? r2_942 : r2_941;
wire r3_472;
assign r3_472 = in[2]? r2_944 : r2_943;
wire r3_473;
assign r3_473 = in[2]? r2_946 : r2_945;
wire r3_474;
assign r3_474 = in[2]? r2_948 : r2_947;
wire r3_475;
assign r3_475 = in[2]? r2_950 : r2_949;
wire r3_476;
assign r3_476 = in[2]? r2_952 : r2_951;
wire r3_477;
assign r3_477 = in[2]? r2_954 : r2_953;
wire r3_478;
assign r3_478 = in[2]? r2_956 : r2_955;
wire r3_479;
assign r3_479 = in[2]? r2_958 : r2_957;
wire r3_480;
assign r3_480 = in[2]? r2_960 : r2_959;
wire r3_481;
assign r3_481 = in[2]? r2_962 : r2_961;
wire r3_482;
assign r3_482 = in[2]? r2_964 : r2_963;
wire r3_483;
assign r3_483 = in[2]? r2_966 : r2_965;
wire r3_484;
assign r3_484 = in[2]? r2_968 : r2_967;
wire r3_485;
assign r3_485 = in[2]? r2_970 : r2_969;
wire r3_486;
assign r3_486 = in[2]? r2_972 : r2_971;
wire r3_487;
assign r3_487 = in[2]? r2_974 : r2_973;
wire r3_488;
assign r3_488 = in[2]? r2_976 : r2_975;
wire r3_489;
assign r3_489 = in[2]? r2_978 : r2_977;
wire r3_490;
assign r3_490 = in[2]? r2_980 : r2_979;
wire r3_491;
assign r3_491 = in[2]? r2_982 : r2_981;
wire r3_492;
assign r3_492 = in[2]? r2_984 : r2_983;
wire r3_493;
assign r3_493 = in[2]? r2_986 : r2_985;
wire r3_494;
assign r3_494 = in[2]? r2_988 : r2_987;
wire r3_495;
assign r3_495 = in[2]? r2_990 : r2_989;
wire r3_496;
assign r3_496 = in[2]? r2_992 : r2_991;
wire r3_497;
assign r3_497 = in[2]? r2_994 : r2_993;
wire r3_498;
assign r3_498 = in[2]? r2_996 : r2_995;
wire r3_499;
assign r3_499 = in[2]? r2_998 : r2_997;
wire r3_500;
assign r3_500 = in[2]? r2_1000 : r2_999;
wire r3_501;
assign r3_501 = in[2]? r2_1002 : r2_1001;
wire r3_502;
assign r3_502 = in[2]? r2_1004 : r2_1003;
wire r3_503;
assign r3_503 = in[2]? r2_1006 : r2_1005;
wire r3_504;
assign r3_504 = in[2]? r2_1008 : r2_1007;
wire r3_505;
assign r3_505 = in[2]? r2_1010 : r2_1009;
wire r3_506;
assign r3_506 = in[2]? r2_1012 : r2_1011;
wire r3_507;
assign r3_507 = in[2]? r2_1014 : r2_1013;
wire r3_508;
assign r3_508 = in[2]? r2_1016 : r2_1015;
wire r3_509;
assign r3_509 = in[2]? r2_1018 : r2_1017;
wire r3_510;
assign r3_510 = in[2]? r2_1020 : r2_1019;
wire r3_511;
assign r3_511 = in[2]? r2_1022 : r2_1021;
wire r3_512;
assign r3_512 = in[2]? r2_1024 : r2_1023;
wire r3_513;
assign r3_513 = in[2]? r2_1026 : r2_1025;
wire r3_514;
assign r3_514 = in[2]? r2_1028 : r2_1027;
wire r3_515;
assign r3_515 = in[2]? r2_1030 : r2_1029;
wire r3_516;
assign r3_516 = in[2]? r2_1032 : r2_1031;
wire r3_517;
assign r3_517 = in[2]? r2_1034 : r2_1033;
wire r3_518;
assign r3_518 = in[2]? r2_1036 : r2_1035;
wire r3_519;
assign r3_519 = in[2]? r2_1038 : r2_1037;
wire r3_520;
assign r3_520 = in[2]? r2_1040 : r2_1039;
wire r3_521;
assign r3_521 = in[2]? r2_1042 : r2_1041;
wire r3_522;
assign r3_522 = in[2]? r2_1044 : r2_1043;
wire r3_523;
assign r3_523 = in[2]? r2_1046 : r2_1045;
wire r3_524;
assign r3_524 = in[2]? r2_1048 : r2_1047;
wire r3_525;
assign r3_525 = in[2]? r2_1050 : r2_1049;
wire r3_526;
assign r3_526 = in[2]? r2_1052 : r2_1051;
wire r3_527;
assign r3_527 = in[2]? r2_1054 : r2_1053;
wire r3_528;
assign r3_528 = in[2]? r2_1056 : r2_1055;
wire r3_529;
assign r3_529 = in[2]? r2_1058 : r2_1057;
wire r3_530;
assign r3_530 = in[2]? r2_1060 : r2_1059;
wire r3_531;
assign r3_531 = in[2]? r2_1062 : r2_1061;
wire r3_532;
assign r3_532 = in[2]? r2_1064 : r2_1063;
wire r3_533;
assign r3_533 = in[2]? r2_1066 : r2_1065;
wire r3_534;
assign r3_534 = in[2]? r2_1068 : r2_1067;
wire r3_535;
assign r3_535 = in[2]? r2_1070 : r2_1069;
wire r3_536;
assign r3_536 = in[2]? r2_1072 : r2_1071;
wire r3_537;
assign r3_537 = in[2]? r2_1074 : r2_1073;
wire r3_538;
assign r3_538 = in[2]? r2_1076 : r2_1075;
wire r3_539;
assign r3_539 = in[2]? r2_1078 : r2_1077;
wire r3_540;
assign r3_540 = in[2]? r2_1080 : r2_1079;
wire r3_541;
assign r3_541 = in[2]? r2_1082 : r2_1081;
wire r3_542;
assign r3_542 = in[2]? r2_1084 : r2_1083;
wire r3_543;
assign r3_543 = in[2]? r2_1086 : r2_1085;
wire r3_544;
assign r3_544 = in[2]? r2_1088 : r2_1087;
wire r3_545;
assign r3_545 = in[2]? r2_1090 : r2_1089;
wire r3_546;
assign r3_546 = in[2]? r2_1092 : r2_1091;
wire r3_547;
assign r3_547 = in[2]? r2_1094 : r2_1093;
wire r3_548;
assign r3_548 = in[2]? r2_1096 : r2_1095;
wire r3_549;
assign r3_549 = in[2]? r2_1098 : r2_1097;
wire r3_550;
assign r3_550 = in[2]? r2_1100 : r2_1099;
wire r3_551;
assign r3_551 = in[2]? r2_1102 : r2_1101;
wire r3_552;
assign r3_552 = in[2]? r2_1104 : r2_1103;
wire r3_553;
assign r3_553 = in[2]? r2_1106 : r2_1105;
wire r3_554;
assign r3_554 = in[2]? r2_1108 : r2_1107;
wire r3_555;
assign r3_555 = in[2]? r2_1110 : r2_1109;
wire r3_556;
assign r3_556 = in[2]? r2_1112 : r2_1111;
wire r3_557;
assign r3_557 = in[2]? r2_1114 : r2_1113;
wire r3_558;
assign r3_558 = in[2]? r2_1116 : r2_1115;
wire r3_559;
assign r3_559 = in[2]? r2_1118 : r2_1117;
wire r3_560;
assign r3_560 = in[2]? r2_1120 : r2_1119;
wire r3_561;
assign r3_561 = in[2]? r2_1122 : r2_1121;
wire r3_562;
assign r3_562 = in[2]? r2_1124 : r2_1123;
wire r3_563;
assign r3_563 = in[2]? r2_1126 : r2_1125;
wire r3_564;
assign r3_564 = in[2]? r2_1128 : r2_1127;
wire r3_565;
assign r3_565 = in[2]? r2_1130 : r2_1129;
wire r3_566;
assign r3_566 = in[2]? r2_1132 : r2_1131;
wire r3_567;
assign r3_567 = in[2]? r2_1134 : r2_1133;
wire r3_568;
assign r3_568 = in[2]? r2_1136 : r2_1135;
wire r3_569;
assign r3_569 = in[2]? r2_1138 : r2_1137;
wire r3_570;
assign r3_570 = in[2]? r2_1140 : r2_1139;
wire r3_571;
assign r3_571 = in[2]? r2_1142 : r2_1141;
wire r3_572;
assign r3_572 = in[2]? r2_1144 : r2_1143;
wire r3_573;
assign r3_573 = in[2]? r2_1146 : r2_1145;
wire r3_574;
assign r3_574 = in[2]? r2_1148 : r2_1147;
wire r3_575;
assign r3_575 = in[2]? r2_1150 : r2_1149;
wire r3_576;
assign r3_576 = in[2]? r2_1152 : r2_1151;
wire r3_577;
assign r3_577 = in[2]? r2_1154 : r2_1153;
wire r3_578;
assign r3_578 = in[2]? r2_1156 : r2_1155;
wire r3_579;
assign r3_579 = in[2]? r2_1158 : r2_1157;
wire r3_580;
assign r3_580 = in[2]? r2_1160 : r2_1159;
wire r3_581;
assign r3_581 = in[2]? r2_1162 : r2_1161;
wire r3_582;
assign r3_582 = in[2]? r2_1164 : r2_1163;
wire r3_583;
assign r3_583 = in[2]? r2_1166 : r2_1165;
wire r3_584;
assign r3_584 = in[2]? r2_1168 : r2_1167;
wire r3_585;
assign r3_585 = in[2]? r2_1170 : r2_1169;
wire r3_586;
assign r3_586 = in[2]? r2_1172 : r2_1171;
wire r3_587;
assign r3_587 = in[2]? r2_1174 : r2_1173;
wire r3_588;
assign r3_588 = in[2]? r2_1176 : r2_1175;
wire r3_589;
assign r3_589 = in[2]? r2_1178 : r2_1177;
wire r3_590;
assign r3_590 = in[2]? r2_1180 : r2_1179;
wire r3_591;
assign r3_591 = in[2]? r2_1182 : r2_1181;
wire r3_592;
assign r3_592 = in[2]? r2_1184 : r2_1183;
wire r3_593;
assign r3_593 = in[2]? r2_1186 : r2_1185;
wire r3_594;
assign r3_594 = in[2]? r2_1188 : r2_1187;
wire r3_595;
assign r3_595 = in[2]? r2_1190 : r2_1189;
wire r3_596;
assign r3_596 = in[2]? r2_1192 : r2_1191;
wire r3_597;
assign r3_597 = in[2]? r2_1194 : r2_1193;
wire r3_598;
assign r3_598 = in[2]? r2_1196 : r2_1195;
wire r3_599;
assign r3_599 = in[2]? r2_1198 : r2_1197;
wire r3_600;
assign r3_600 = in[2]? r2_1200 : r2_1199;
wire r3_601;
assign r3_601 = in[2]? r2_1202 : r2_1201;
wire r3_602;
assign r3_602 = in[2]? r2_1204 : r2_1203;
wire r3_603;
assign r3_603 = in[2]? r2_1206 : r2_1205;
wire r3_604;
assign r3_604 = in[2]? r2_1208 : r2_1207;
wire r3_605;
assign r3_605 = in[2]? r2_1210 : r2_1209;
wire r3_606;
assign r3_606 = in[2]? r2_1212 : r2_1211;
wire r3_607;
assign r3_607 = in[2]? r2_1214 : r2_1213;
wire r3_608;
assign r3_608 = in[2]? r2_1216 : r2_1215;
wire r3_609;
assign r3_609 = in[2]? r2_1218 : r2_1217;
wire r3_610;
assign r3_610 = in[2]? r2_1220 : r2_1219;
wire r3_611;
assign r3_611 = in[2]? r2_1222 : r2_1221;
wire r3_612;
assign r3_612 = in[2]? r2_1224 : r2_1223;
wire r3_613;
assign r3_613 = in[2]? r2_1226 : r2_1225;
wire r3_614;
assign r3_614 = in[2]? r2_1228 : r2_1227;
wire r3_615;
assign r3_615 = in[2]? r2_1230 : r2_1229;
wire r3_616;
assign r3_616 = in[2]? r2_1232 : r2_1231;
wire r3_617;
assign r3_617 = in[2]? r2_1234 : r2_1233;
wire r3_618;
assign r3_618 = in[2]? r2_1236 : r2_1235;
wire r3_619;
assign r3_619 = in[2]? r2_1238 : r2_1237;
wire r3_620;
assign r3_620 = in[2]? r2_1240 : r2_1239;
wire r3_621;
assign r3_621 = in[2]? r2_1242 : r2_1241;
wire r3_622;
assign r3_622 = in[2]? r2_1244 : r2_1243;
wire r3_623;
assign r3_623 = in[2]? r2_1246 : r2_1245;
wire r3_624;
assign r3_624 = in[2]? r2_1248 : r2_1247;
wire r3_625;
assign r3_625 = in[2]? r2_1250 : r2_1249;
wire r3_626;
assign r3_626 = in[2]? r2_1252 : r2_1251;
wire r3_627;
assign r3_627 = in[2]? r2_1254 : r2_1253;
wire r3_628;
assign r3_628 = in[2]? r2_1256 : r2_1255;
wire r3_629;
assign r3_629 = in[2]? r2_1258 : r2_1257;
wire r3_630;
assign r3_630 = in[2]? r2_1260 : r2_1259;
wire r3_631;
assign r3_631 = in[2]? r2_1262 : r2_1261;
wire r3_632;
assign r3_632 = in[2]? r2_1264 : r2_1263;
wire r3_633;
assign r3_633 = in[2]? r2_1266 : r2_1265;
wire r3_634;
assign r3_634 = in[2]? r2_1268 : r2_1267;
wire r3_635;
assign r3_635 = in[2]? r2_1270 : r2_1269;
wire r3_636;
assign r3_636 = in[2]? r2_1272 : r2_1271;
wire r3_637;
assign r3_637 = in[2]? r2_1274 : r2_1273;
wire r3_638;
assign r3_638 = in[2]? r2_1276 : r2_1275;
wire r3_639;
assign r3_639 = in[2]? r2_1278 : r2_1277;
wire r3_640;
assign r3_640 = in[2]? r2_1280 : r2_1279;
wire r3_641;
assign r3_641 = in[2]? r2_1282 : r2_1281;
wire r3_642;
assign r3_642 = in[2]? r2_1284 : r2_1283;
wire r3_643;
assign r3_643 = in[2]? r2_1286 : r2_1285;
wire r3_644;
assign r3_644 = in[2]? r2_1288 : r2_1287;
wire r3_645;
assign r3_645 = in[2]? r2_1290 : r2_1289;
wire r3_646;
assign r3_646 = in[2]? r2_1292 : r2_1291;
wire r3_647;
assign r3_647 = in[2]? r2_1294 : r2_1293;
wire r3_648;
assign r3_648 = in[2]? r2_1296 : r2_1295;
wire r3_649;
assign r3_649 = in[2]? r2_1298 : r2_1297;
wire r3_650;
assign r3_650 = in[2]? r2_1300 : r2_1299;
wire r3_651;
assign r3_651 = in[2]? r2_1302 : r2_1301;
wire r3_652;
assign r3_652 = in[2]? r2_1304 : r2_1303;
wire r3_653;
assign r3_653 = in[2]? r2_1306 : r2_1305;
wire r3_654;
assign r3_654 = in[2]? r2_1308 : r2_1307;
wire r3_655;
assign r3_655 = in[2]? r2_1310 : r2_1309;
wire r3_656;
assign r3_656 = in[2]? r2_1312 : r2_1311;
wire r3_657;
assign r3_657 = in[2]? r2_1314 : r2_1313;
wire r3_658;
assign r3_658 = in[2]? r2_1316 : r2_1315;
wire r3_659;
assign r3_659 = in[2]? r2_1318 : r2_1317;
wire r3_660;
assign r3_660 = in[2]? r2_1320 : r2_1319;
wire r3_661;
assign r3_661 = in[2]? r2_1322 : r2_1321;
wire r3_662;
assign r3_662 = in[2]? r2_1324 : r2_1323;
wire r3_663;
assign r3_663 = in[2]? r2_1326 : r2_1325;
wire r3_664;
assign r3_664 = in[2]? r2_1328 : r2_1327;
wire r3_665;
assign r3_665 = in[2]? r2_1330 : r2_1329;
wire r3_666;
assign r3_666 = in[2]? r2_1332 : r2_1331;
wire r3_667;
assign r3_667 = in[2]? r2_1334 : r2_1333;
wire r3_668;
assign r3_668 = in[2]? r2_1336 : r2_1335;
wire r3_669;
assign r3_669 = in[2]? r2_1338 : r2_1337;
wire r3_670;
assign r3_670 = in[2]? r2_1340 : r2_1339;
wire r3_671;
assign r3_671 = in[2]? r2_1342 : r2_1341;
wire r3_672;
assign r3_672 = in[2]? r2_1344 : r2_1343;
wire r3_673;
assign r3_673 = in[2]? r2_1346 : r2_1345;
wire r3_674;
assign r3_674 = in[2]? r2_1348 : r2_1347;
wire r3_675;
assign r3_675 = in[2]? r2_1350 : r2_1349;
wire r3_676;
assign r3_676 = in[2]? r2_1352 : r2_1351;
wire r3_677;
assign r3_677 = in[2]? r2_1354 : r2_1353;
wire r3_678;
assign r3_678 = in[2]? r2_1356 : r2_1355;
wire r3_679;
assign r3_679 = in[2]? r2_1358 : r2_1357;
wire r3_680;
assign r3_680 = in[2]? r2_1360 : r2_1359;
wire r3_681;
assign r3_681 = in[2]? r2_1362 : r2_1361;
wire r3_682;
assign r3_682 = in[2]? r2_1364 : r2_1363;
wire r3_683;
assign r3_683 = in[2]? r2_1366 : r2_1365;
wire r3_684;
assign r3_684 = in[2]? r2_1368 : r2_1367;
wire r3_685;
assign r3_685 = in[2]? r2_1370 : r2_1369;
wire r3_686;
assign r3_686 = in[2]? r2_1372 : r2_1371;
wire r3_687;
assign r3_687 = in[2]? r2_1374 : r2_1373;
wire r3_688;
assign r3_688 = in[2]? r2_1376 : r2_1375;
wire r3_689;
assign r3_689 = in[2]? r2_1378 : r2_1377;
wire r3_690;
assign r3_690 = in[2]? r2_1380 : r2_1379;
wire r3_691;
assign r3_691 = in[2]? r2_1382 : r2_1381;
wire r3_692;
assign r3_692 = in[2]? r2_1384 : r2_1383;
wire r3_693;
assign r3_693 = in[2]? r2_1386 : r2_1385;
wire r3_694;
assign r3_694 = in[2]? r2_1388 : r2_1387;
wire r3_695;
assign r3_695 = in[2]? r2_1390 : r2_1389;
wire r3_696;
assign r3_696 = in[2]? r2_1392 : r2_1391;
wire r3_697;
assign r3_697 = in[2]? r2_1394 : r2_1393;
wire r3_698;
assign r3_698 = in[2]? r2_1396 : r2_1395;
wire r3_699;
assign r3_699 = in[2]? r2_1398 : r2_1397;
wire r3_700;
assign r3_700 = in[2]? r2_1400 : r2_1399;
wire r3_701;
assign r3_701 = in[2]? r2_1402 : r2_1401;
wire r3_702;
assign r3_702 = in[2]? r2_1404 : r2_1403;
wire r3_703;
assign r3_703 = in[2]? r2_1406 : r2_1405;
wire r3_704;
assign r3_704 = in[2]? r2_1408 : r2_1407;
wire r3_705;
assign r3_705 = in[2]? r2_1410 : r2_1409;
wire r3_706;
assign r3_706 = in[2]? r2_1412 : r2_1411;
wire r3_707;
assign r3_707 = in[2]? r2_1414 : r2_1413;
wire r3_708;
assign r3_708 = in[2]? r2_1416 : r2_1415;
wire r3_709;
assign r3_709 = in[2]? r2_1418 : r2_1417;
wire r3_710;
assign r3_710 = in[2]? r2_1420 : r2_1419;
wire r3_711;
assign r3_711 = in[2]? r2_1422 : r2_1421;
wire r3_712;
assign r3_712 = in[2]? r2_1424 : r2_1423;
wire r3_713;
assign r3_713 = in[2]? r2_1426 : r2_1425;
wire r3_714;
assign r3_714 = in[2]? r2_1428 : r2_1427;
wire r3_715;
assign r3_715 = in[2]? r2_1430 : r2_1429;
wire r3_716;
assign r3_716 = in[2]? r2_1432 : r2_1431;
wire r3_717;
assign r3_717 = in[2]? r2_1434 : r2_1433;
wire r3_718;
assign r3_718 = in[2]? r2_1436 : r2_1435;
wire r3_719;
assign r3_719 = in[2]? r2_1438 : r2_1437;
wire r3_720;
assign r3_720 = in[2]? r2_1440 : r2_1439;
wire r3_721;
assign r3_721 = in[2]? r2_1442 : r2_1441;
wire r3_722;
assign r3_722 = in[2]? r2_1444 : r2_1443;
wire r3_723;
assign r3_723 = in[2]? r2_1446 : r2_1445;
wire r3_724;
assign r3_724 = in[2]? r2_1448 : r2_1447;
wire r3_725;
assign r3_725 = in[2]? r2_1450 : r2_1449;
wire r3_726;
assign r3_726 = in[2]? r2_1452 : r2_1451;
wire r3_727;
assign r3_727 = in[2]? r2_1454 : r2_1453;
wire r3_728;
assign r3_728 = in[2]? r2_1456 : r2_1455;
wire r3_729;
assign r3_729 = in[2]? r2_1458 : r2_1457;
wire r3_730;
assign r3_730 = in[2]? r2_1460 : r2_1459;
wire r3_731;
assign r3_731 = in[2]? r2_1462 : r2_1461;
wire r3_732;
assign r3_732 = in[2]? r2_1464 : r2_1463;
wire r3_733;
assign r3_733 = in[2]? r2_1466 : r2_1465;
wire r3_734;
assign r3_734 = in[2]? r2_1468 : r2_1467;
wire r3_735;
assign r3_735 = in[2]? r2_1470 : r2_1469;
wire r3_736;
assign r3_736 = in[2]? r2_1472 : r2_1471;
wire r3_737;
assign r3_737 = in[2]? r2_1474 : r2_1473;
wire r3_738;
assign r3_738 = in[2]? r2_1476 : r2_1475;
wire r3_739;
assign r3_739 = in[2]? r2_1478 : r2_1477;
wire r3_740;
assign r3_740 = in[2]? r2_1480 : r2_1479;
wire r3_741;
assign r3_741 = in[2]? r2_1482 : r2_1481;
wire r3_742;
assign r3_742 = in[2]? r2_1484 : r2_1483;
wire r3_743;
assign r3_743 = in[2]? r2_1486 : r2_1485;
wire r3_744;
assign r3_744 = in[2]? r2_1488 : r2_1487;
wire r3_745;
assign r3_745 = in[2]? r2_1490 : r2_1489;
wire r3_746;
assign r3_746 = in[2]? r2_1492 : r2_1491;
wire r3_747;
assign r3_747 = in[2]? r2_1494 : r2_1493;
wire r3_748;
assign r3_748 = in[2]? r2_1496 : r2_1495;
wire r3_749;
assign r3_749 = in[2]? r2_1498 : r2_1497;
wire r3_750;
assign r3_750 = in[2]? r2_1500 : r2_1499;
wire r3_751;
assign r3_751 = in[2]? r2_1502 : r2_1501;
wire r3_752;
assign r3_752 = in[2]? r2_1504 : r2_1503;
wire r3_753;
assign r3_753 = in[2]? r2_1506 : r2_1505;
wire r3_754;
assign r3_754 = in[2]? r2_1508 : r2_1507;
wire r3_755;
assign r3_755 = in[2]? r2_1510 : r2_1509;
wire r3_756;
assign r3_756 = in[2]? r2_1512 : r2_1511;
wire r3_757;
assign r3_757 = in[2]? r2_1514 : r2_1513;
wire r3_758;
assign r3_758 = in[2]? r2_1516 : r2_1515;
wire r3_759;
assign r3_759 = in[2]? r2_1518 : r2_1517;
wire r3_760;
assign r3_760 = in[2]? r2_1520 : r2_1519;
wire r3_761;
assign r3_761 = in[2]? r2_1522 : r2_1521;
wire r3_762;
assign r3_762 = in[2]? r2_1524 : r2_1523;
wire r3_763;
assign r3_763 = in[2]? r2_1526 : r2_1525;
wire r3_764;
assign r3_764 = in[2]? r2_1528 : r2_1527;
wire r3_765;
assign r3_765 = in[2]? r2_1530 : r2_1529;
wire r3_766;
assign r3_766 = in[2]? r2_1532 : r2_1531;
wire r3_767;
assign r3_767 = in[2]? r2_1534 : r2_1533;
wire r3_768;
assign r3_768 = in[2]? r2_1536 : r2_1535;
wire r3_769;
assign r3_769 = in[2]? r2_1538 : r2_1537;
wire r3_770;
assign r3_770 = in[2]? r2_1540 : r2_1539;
wire r3_771;
assign r3_771 = in[2]? r2_1542 : r2_1541;
wire r3_772;
assign r3_772 = in[2]? r2_1544 : r2_1543;
wire r3_773;
assign r3_773 = in[2]? r2_1546 : r2_1545;
wire r3_774;
assign r3_774 = in[2]? r2_1548 : r2_1547;
wire r3_775;
assign r3_775 = in[2]? r2_1550 : r2_1549;
wire r3_776;
assign r3_776 = in[2]? r2_1552 : r2_1551;
wire r3_777;
assign r3_777 = in[2]? r2_1554 : r2_1553;
wire r3_778;
assign r3_778 = in[2]? r2_1556 : r2_1555;
wire r3_779;
assign r3_779 = in[2]? r2_1558 : r2_1557;
wire r3_780;
assign r3_780 = in[2]? r2_1560 : r2_1559;
wire r3_781;
assign r3_781 = in[2]? r2_1562 : r2_1561;
wire r3_782;
assign r3_782 = in[2]? r2_1564 : r2_1563;
wire r3_783;
assign r3_783 = in[2]? r2_1566 : r2_1565;
wire r3_784;
assign r3_784 = in[2]? r2_1568 : r2_1567;
wire r3_785;
assign r3_785 = in[2]? r2_1570 : r2_1569;
wire r3_786;
assign r3_786 = in[2]? r2_1572 : r2_1571;
wire r3_787;
assign r3_787 = in[2]? r2_1574 : r2_1573;
wire r3_788;
assign r3_788 = in[2]? r2_1576 : r2_1575;
wire r3_789;
assign r3_789 = in[2]? r2_1578 : r2_1577;
wire r3_790;
assign r3_790 = in[2]? r2_1580 : r2_1579;
wire r3_791;
assign r3_791 = in[2]? r2_1582 : r2_1581;
wire r3_792;
assign r3_792 = in[2]? r2_1584 : r2_1583;
wire r3_793;
assign r3_793 = in[2]? r2_1586 : r2_1585;
wire r3_794;
assign r3_794 = in[2]? r2_1588 : r2_1587;
wire r3_795;
assign r3_795 = in[2]? r2_1590 : r2_1589;
wire r3_796;
assign r3_796 = in[2]? r2_1592 : r2_1591;
wire r3_797;
assign r3_797 = in[2]? r2_1594 : r2_1593;
wire r3_798;
assign r3_798 = in[2]? r2_1596 : r2_1595;
wire r3_799;
assign r3_799 = in[2]? r2_1598 : r2_1597;
wire r3_800;
assign r3_800 = in[2]? r2_1600 : r2_1599;
wire r3_801;
assign r3_801 = in[2]? r2_1602 : r2_1601;
wire r3_802;
assign r3_802 = in[2]? r2_1604 : r2_1603;
wire r3_803;
assign r3_803 = in[2]? r2_1606 : r2_1605;
wire r3_804;
assign r3_804 = in[2]? r2_1608 : r2_1607;
wire r3_805;
assign r3_805 = in[2]? r2_1610 : r2_1609;
wire r3_806;
assign r3_806 = in[2]? r2_1612 : r2_1611;
wire r3_807;
assign r3_807 = in[2]? r2_1614 : r2_1613;
wire r3_808;
assign r3_808 = in[2]? r2_1616 : r2_1615;
wire r3_809;
assign r3_809 = in[2]? r2_1618 : r2_1617;
wire r3_810;
assign r3_810 = in[2]? r2_1620 : r2_1619;
wire r3_811;
assign r3_811 = in[2]? r2_1622 : r2_1621;
wire r3_812;
assign r3_812 = in[2]? r2_1624 : r2_1623;
wire r3_813;
assign r3_813 = in[2]? r2_1626 : r2_1625;
wire r3_814;
assign r3_814 = in[2]? r2_1628 : r2_1627;
wire r3_815;
assign r3_815 = in[2]? r2_1630 : r2_1629;
wire r3_816;
assign r3_816 = in[2]? r2_1632 : r2_1631;
wire r3_817;
assign r3_817 = in[2]? r2_1634 : r2_1633;
wire r3_818;
assign r3_818 = in[2]? r2_1636 : r2_1635;
wire r3_819;
assign r3_819 = in[2]? r2_1638 : r2_1637;
wire r3_820;
assign r3_820 = in[2]? r2_1640 : r2_1639;
wire r3_821;
assign r3_821 = in[2]? r2_1642 : r2_1641;
wire r3_822;
assign r3_822 = in[2]? r2_1644 : r2_1643;
wire r3_823;
assign r3_823 = in[2]? r2_1646 : r2_1645;
wire r3_824;
assign r3_824 = in[2]? r2_1648 : r2_1647;
wire r3_825;
assign r3_825 = in[2]? r2_1650 : r2_1649;
wire r3_826;
assign r3_826 = in[2]? r2_1652 : r2_1651;
wire r3_827;
assign r3_827 = in[2]? r2_1654 : r2_1653;
wire r3_828;
assign r3_828 = in[2]? r2_1656 : r2_1655;
wire r3_829;
assign r3_829 = in[2]? r2_1658 : r2_1657;
wire r3_830;
assign r3_830 = in[2]? r2_1660 : r2_1659;
wire r3_831;
assign r3_831 = in[2]? r2_1662 : r2_1661;
wire r3_832;
assign r3_832 = in[2]? r2_1664 : r2_1663;
wire r3_833;
assign r3_833 = in[2]? r2_1666 : r2_1665;
wire r3_834;
assign r3_834 = in[2]? r2_1668 : r2_1667;
wire r3_835;
assign r3_835 = in[2]? r2_1670 : r2_1669;
wire r3_836;
assign r3_836 = in[2]? r2_1672 : r2_1671;
wire r3_837;
assign r3_837 = in[2]? r2_1674 : r2_1673;
wire r3_838;
assign r3_838 = in[2]? r2_1676 : r2_1675;
wire r3_839;
assign r3_839 = in[2]? r2_1678 : r2_1677;
wire r3_840;
assign r3_840 = in[2]? r2_1680 : r2_1679;
wire r3_841;
assign r3_841 = in[2]? r2_1682 : r2_1681;
wire r3_842;
assign r3_842 = in[2]? r2_1684 : r2_1683;
wire r3_843;
assign r3_843 = in[2]? r2_1686 : r2_1685;
wire r3_844;
assign r3_844 = in[2]? r2_1688 : r2_1687;
wire r3_845;
assign r3_845 = in[2]? r2_1690 : r2_1689;
wire r3_846;
assign r3_846 = in[2]? r2_1692 : r2_1691;
wire r3_847;
assign r3_847 = in[2]? r2_1694 : r2_1693;
wire r3_848;
assign r3_848 = in[2]? r2_1696 : r2_1695;
wire r3_849;
assign r3_849 = in[2]? r2_1698 : r2_1697;
wire r3_850;
assign r3_850 = in[2]? r2_1700 : r2_1699;
wire r3_851;
assign r3_851 = in[2]? r2_1702 : r2_1701;
wire r3_852;
assign r3_852 = in[2]? r2_1704 : r2_1703;
wire r3_853;
assign r3_853 = in[2]? r2_1706 : r2_1705;
wire r3_854;
assign r3_854 = in[2]? r2_1708 : r2_1707;
wire r3_855;
assign r3_855 = in[2]? r2_1710 : r2_1709;
wire r3_856;
assign r3_856 = in[2]? r2_1712 : r2_1711;
wire r3_857;
assign r3_857 = in[2]? r2_1714 : r2_1713;
wire r3_858;
assign r3_858 = in[2]? r2_1716 : r2_1715;
wire r3_859;
assign r3_859 = in[2]? r2_1718 : r2_1717;
wire r3_860;
assign r3_860 = in[2]? r2_1720 : r2_1719;
wire r3_861;
assign r3_861 = in[2]? r2_1722 : r2_1721;
wire r3_862;
assign r3_862 = in[2]? r2_1724 : r2_1723;
wire r3_863;
assign r3_863 = in[2]? r2_1726 : r2_1725;
wire r3_864;
assign r3_864 = in[2]? r2_1728 : r2_1727;
wire r3_865;
assign r3_865 = in[2]? r2_1730 : r2_1729;
wire r3_866;
assign r3_866 = in[2]? r2_1732 : r2_1731;
wire r3_867;
assign r3_867 = in[2]? r2_1734 : r2_1733;
wire r3_868;
assign r3_868 = in[2]? r2_1736 : r2_1735;
wire r3_869;
assign r3_869 = in[2]? r2_1738 : r2_1737;
wire r3_870;
assign r3_870 = in[2]? r2_1740 : r2_1739;
wire r3_871;
assign r3_871 = in[2]? r2_1742 : r2_1741;
wire r3_872;
assign r3_872 = in[2]? r2_1744 : r2_1743;
wire r3_873;
assign r3_873 = in[2]? r2_1746 : r2_1745;
wire r3_874;
assign r3_874 = in[2]? r2_1748 : r2_1747;
wire r3_875;
assign r3_875 = in[2]? r2_1750 : r2_1749;
wire r3_876;
assign r3_876 = in[2]? r2_1752 : r2_1751;
wire r3_877;
assign r3_877 = in[2]? r2_1754 : r2_1753;
wire r3_878;
assign r3_878 = in[2]? r2_1756 : r2_1755;
wire r3_879;
assign r3_879 = in[2]? r2_1758 : r2_1757;
wire r3_880;
assign r3_880 = in[2]? r2_1760 : r2_1759;
wire r3_881;
assign r3_881 = in[2]? r2_1762 : r2_1761;
wire r3_882;
assign r3_882 = in[2]? r2_1764 : r2_1763;
wire r3_883;
assign r3_883 = in[2]? r2_1766 : r2_1765;
wire r3_884;
assign r3_884 = in[2]? r2_1768 : r2_1767;
wire r3_885;
assign r3_885 = in[2]? r2_1770 : r2_1769;
wire r3_886;
assign r3_886 = in[2]? r2_1772 : r2_1771;
wire r3_887;
assign r3_887 = in[2]? r2_1774 : r2_1773;
wire r3_888;
assign r3_888 = in[2]? r2_1776 : r2_1775;
wire r3_889;
assign r3_889 = in[2]? r2_1778 : r2_1777;
wire r3_890;
assign r3_890 = in[2]? r2_1780 : r2_1779;
wire r3_891;
assign r3_891 = in[2]? r2_1782 : r2_1781;
wire r3_892;
assign r3_892 = in[2]? r2_1784 : r2_1783;
wire r3_893;
assign r3_893 = in[2]? r2_1786 : r2_1785;
wire r3_894;
assign r3_894 = in[2]? r2_1788 : r2_1787;
wire r3_895;
assign r3_895 = in[2]? r2_1790 : r2_1789;
wire r3_896;
assign r3_896 = in[2]? r2_1792 : r2_1791;
wire r3_897;
assign r3_897 = in[2]? r2_1794 : r2_1793;
wire r3_898;
assign r3_898 = in[2]? r2_1796 : r2_1795;
wire r3_899;
assign r3_899 = in[2]? r2_1798 : r2_1797;
wire r3_900;
assign r3_900 = in[2]? r2_1800 : r2_1799;
wire r3_901;
assign r3_901 = in[2]? r2_1802 : r2_1801;
wire r3_902;
assign r3_902 = in[2]? r2_1804 : r2_1803;
wire r3_903;
assign r3_903 = in[2]? r2_1806 : r2_1805;
wire r3_904;
assign r3_904 = in[2]? r2_1808 : r2_1807;
wire r3_905;
assign r3_905 = in[2]? r2_1810 : r2_1809;
wire r3_906;
assign r3_906 = in[2]? r2_1812 : r2_1811;
wire r3_907;
assign r3_907 = in[2]? r2_1814 : r2_1813;
wire r3_908;
assign r3_908 = in[2]? r2_1816 : r2_1815;
wire r3_909;
assign r3_909 = in[2]? r2_1818 : r2_1817;
wire r3_910;
assign r3_910 = in[2]? r2_1820 : r2_1819;
wire r3_911;
assign r3_911 = in[2]? r2_1822 : r2_1821;
wire r3_912;
assign r3_912 = in[2]? r2_1824 : r2_1823;
wire r3_913;
assign r3_913 = in[2]? r2_1826 : r2_1825;
wire r3_914;
assign r3_914 = in[2]? r2_1828 : r2_1827;
wire r3_915;
assign r3_915 = in[2]? r2_1830 : r2_1829;
wire r3_916;
assign r3_916 = in[2]? r2_1832 : r2_1831;
wire r3_917;
assign r3_917 = in[2]? r2_1834 : r2_1833;
wire r3_918;
assign r3_918 = in[2]? r2_1836 : r2_1835;
wire r3_919;
assign r3_919 = in[2]? r2_1838 : r2_1837;
wire r3_920;
assign r3_920 = in[2]? r2_1840 : r2_1839;
wire r3_921;
assign r3_921 = in[2]? r2_1842 : r2_1841;
wire r3_922;
assign r3_922 = in[2]? r2_1844 : r2_1843;
wire r3_923;
assign r3_923 = in[2]? r2_1846 : r2_1845;
wire r3_924;
assign r3_924 = in[2]? r2_1848 : r2_1847;
wire r3_925;
assign r3_925 = in[2]? r2_1850 : r2_1849;
wire r3_926;
assign r3_926 = in[2]? r2_1852 : r2_1851;
wire r3_927;
assign r3_927 = in[2]? r2_1854 : r2_1853;
wire r3_928;
assign r3_928 = in[2]? r2_1856 : r2_1855;
wire r3_929;
assign r3_929 = in[2]? r2_1858 : r2_1857;
wire r3_930;
assign r3_930 = in[2]? r2_1860 : r2_1859;
wire r3_931;
assign r3_931 = in[2]? r2_1862 : r2_1861;
wire r3_932;
assign r3_932 = in[2]? r2_1864 : r2_1863;
wire r3_933;
assign r3_933 = in[2]? r2_1866 : r2_1865;
wire r3_934;
assign r3_934 = in[2]? r2_1868 : r2_1867;
wire r3_935;
assign r3_935 = in[2]? r2_1870 : r2_1869;
wire r3_936;
assign r3_936 = in[2]? r2_1872 : r2_1871;
wire r3_937;
assign r3_937 = in[2]? r2_1874 : r2_1873;
wire r3_938;
assign r3_938 = in[2]? r2_1876 : r2_1875;
wire r3_939;
assign r3_939 = in[2]? r2_1878 : r2_1877;
wire r3_940;
assign r3_940 = in[2]? r2_1880 : r2_1879;
wire r3_941;
assign r3_941 = in[2]? r2_1882 : r2_1881;
wire r3_942;
assign r3_942 = in[2]? r2_1884 : r2_1883;
wire r3_943;
assign r3_943 = in[2]? r2_1886 : r2_1885;
wire r3_944;
assign r3_944 = in[2]? r2_1888 : r2_1887;
wire r3_945;
assign r3_945 = in[2]? r2_1890 : r2_1889;
wire r3_946;
assign r3_946 = in[2]? r2_1892 : r2_1891;
wire r3_947;
assign r3_947 = in[2]? r2_1894 : r2_1893;
wire r3_948;
assign r3_948 = in[2]? r2_1896 : r2_1895;
wire r3_949;
assign r3_949 = in[2]? r2_1898 : r2_1897;
wire r3_950;
assign r3_950 = in[2]? r2_1900 : r2_1899;
wire r3_951;
assign r3_951 = in[2]? r2_1902 : r2_1901;
wire r3_952;
assign r3_952 = in[2]? r2_1904 : r2_1903;
wire r3_953;
assign r3_953 = in[2]? r2_1906 : r2_1905;
wire r3_954;
assign r3_954 = in[2]? r2_1908 : r2_1907;
wire r3_955;
assign r3_955 = in[2]? r2_1910 : r2_1909;
wire r3_956;
assign r3_956 = in[2]? r2_1912 : r2_1911;
wire r3_957;
assign r3_957 = in[2]? r2_1914 : r2_1913;
wire r3_958;
assign r3_958 = in[2]? r2_1916 : r2_1915;
wire r3_959;
assign r3_959 = in[2]? r2_1918 : r2_1917;
wire r3_960;
assign r3_960 = in[2]? r2_1920 : r2_1919;
wire r3_961;
assign r3_961 = in[2]? r2_1922 : r2_1921;
wire r3_962;
assign r3_962 = in[2]? r2_1924 : r2_1923;
wire r3_963;
assign r3_963 = in[2]? r2_1926 : r2_1925;
wire r3_964;
assign r3_964 = in[2]? r2_1928 : r2_1927;
wire r3_965;
assign r3_965 = in[2]? r2_1930 : r2_1929;
wire r3_966;
assign r3_966 = in[2]? r2_1932 : r2_1931;
wire r3_967;
assign r3_967 = in[2]? r2_1934 : r2_1933;
wire r3_968;
assign r3_968 = in[2]? r2_1936 : r2_1935;
wire r3_969;
assign r3_969 = in[2]? r2_1938 : r2_1937;
wire r3_970;
assign r3_970 = in[2]? r2_1940 : r2_1939;
wire r3_971;
assign r3_971 = in[2]? r2_1942 : r2_1941;
wire r3_972;
assign r3_972 = in[2]? r2_1944 : r2_1943;
wire r3_973;
assign r3_973 = in[2]? r2_1946 : r2_1945;
wire r3_974;
assign r3_974 = in[2]? r2_1948 : r2_1947;
wire r3_975;
assign r3_975 = in[2]? r2_1950 : r2_1949;
wire r3_976;
assign r3_976 = in[2]? r2_1952 : r2_1951;
wire r3_977;
assign r3_977 = in[2]? r2_1954 : r2_1953;
wire r3_978;
assign r3_978 = in[2]? r2_1956 : r2_1955;
wire r3_979;
assign r3_979 = in[2]? r2_1958 : r2_1957;
wire r3_980;
assign r3_980 = in[2]? r2_1960 : r2_1959;
wire r3_981;
assign r3_981 = in[2]? r2_1962 : r2_1961;
wire r3_982;
assign r3_982 = in[2]? r2_1964 : r2_1963;
wire r3_983;
assign r3_983 = in[2]? r2_1966 : r2_1965;
wire r3_984;
assign r3_984 = in[2]? r2_1968 : r2_1967;
wire r3_985;
assign r3_985 = in[2]? r2_1970 : r2_1969;
wire r3_986;
assign r3_986 = in[2]? r2_1972 : r2_1971;
wire r3_987;
assign r3_987 = in[2]? r2_1974 : r2_1973;
wire r3_988;
assign r3_988 = in[2]? r2_1976 : r2_1975;
wire r3_989;
assign r3_989 = in[2]? r2_1978 : r2_1977;
wire r3_990;
assign r3_990 = in[2]? r2_1980 : r2_1979;
wire r3_991;
assign r3_991 = in[2]? r2_1982 : r2_1981;
wire r3_992;
assign r3_992 = in[2]? r2_1984 : r2_1983;
wire r3_993;
assign r3_993 = in[2]? r2_1986 : r2_1985;
wire r3_994;
assign r3_994 = in[2]? r2_1988 : r2_1987;
wire r3_995;
assign r3_995 = in[2]? r2_1990 : r2_1989;
wire r3_996;
assign r3_996 = in[2]? r2_1992 : r2_1991;
wire r3_997;
assign r3_997 = in[2]? r2_1994 : r2_1993;
wire r3_998;
assign r3_998 = in[2]? r2_1996 : r2_1995;
wire r3_999;
assign r3_999 = in[2]? r2_1998 : r2_1997;
wire r3_1000;
assign r3_1000 = in[2]? r2_2000 : r2_1999;
wire r3_1001;
assign r3_1001 = in[2]? r2_2002 : r2_2001;
wire r3_1002;
assign r3_1002 = in[2]? r2_2004 : r2_2003;
wire r3_1003;
assign r3_1003 = in[2]? r2_2006 : r2_2005;
wire r3_1004;
assign r3_1004 = in[2]? r2_2008 : r2_2007;
wire r3_1005;
assign r3_1005 = in[2]? r2_2010 : r2_2009;
wire r3_1006;
assign r3_1006 = in[2]? r2_2012 : r2_2011;
wire r3_1007;
assign r3_1007 = in[2]? r2_2014 : r2_2013;
wire r3_1008;
assign r3_1008 = in[2]? r2_2016 : r2_2015;
wire r3_1009;
assign r3_1009 = in[2]? r2_2018 : r2_2017;
wire r3_1010;
assign r3_1010 = in[2]? r2_2020 : r2_2019;
wire r3_1011;
assign r3_1011 = in[2]? r2_2022 : r2_2021;
wire r3_1012;
assign r3_1012 = in[2]? r2_2024 : r2_2023;
wire r3_1013;
assign r3_1013 = in[2]? r2_2026 : r2_2025;
wire r3_1014;
assign r3_1014 = in[2]? r2_2028 : r2_2027;
wire r3_1015;
assign r3_1015 = in[2]? r2_2030 : r2_2029;
wire r3_1016;
assign r3_1016 = in[2]? r2_2032 : r2_2031;
wire r3_1017;
assign r3_1017 = in[2]? r2_2034 : r2_2033;
wire r3_1018;
assign r3_1018 = in[2]? r2_2036 : r2_2035;
wire r3_1019;
assign r3_1019 = in[2]? r2_2038 : r2_2037;
wire r3_1020;
assign r3_1020 = in[2]? r2_2040 : r2_2039;
wire r3_1021;
assign r3_1021 = in[2]? r2_2042 : r2_2041;
wire r3_1022;
assign r3_1022 = in[2]? r2_2044 : r2_2043;
wire r3_1023;
assign r3_1023 = in[2]? r2_2046 : r2_2045;
wire r3_1024;
assign r3_1024 = in[2]? r2_2048 : r2_2047;
wire r3_1025;
assign r3_1025 = in[2]? r2_2050 : r2_2049;
wire r3_1026;
assign r3_1026 = in[2]? r2_2052 : r2_2051;
wire r3_1027;
assign r3_1027 = in[2]? r2_2054 : r2_2053;
wire r3_1028;
assign r3_1028 = in[2]? r2_2056 : r2_2055;
wire r3_1029;
assign r3_1029 = in[2]? r2_2058 : r2_2057;
wire r3_1030;
assign r3_1030 = in[2]? r2_2060 : r2_2059;
wire r3_1031;
assign r3_1031 = in[2]? r2_2062 : r2_2061;
wire r3_1032;
assign r3_1032 = in[2]? r2_2064 : r2_2063;
wire r3_1033;
assign r3_1033 = in[2]? r2_2066 : r2_2065;
wire r3_1034;
assign r3_1034 = in[2]? r2_2068 : r2_2067;
wire r3_1035;
assign r3_1035 = in[2]? r2_2070 : r2_2069;
wire r3_1036;
assign r3_1036 = in[2]? r2_2072 : r2_2071;
wire r3_1037;
assign r3_1037 = in[2]? r2_2074 : r2_2073;
wire r3_1038;
assign r3_1038 = in[2]? r2_2076 : r2_2075;
wire r3_1039;
assign r3_1039 = in[2]? r2_2078 : r2_2077;
wire r3_1040;
assign r3_1040 = in[2]? r2_2080 : r2_2079;
wire r3_1041;
assign r3_1041 = in[2]? r2_2082 : r2_2081;
wire r3_1042;
assign r3_1042 = in[2]? r2_2084 : r2_2083;
wire r3_1043;
assign r3_1043 = in[2]? r2_2086 : r2_2085;
wire r3_1044;
assign r3_1044 = in[2]? r2_2088 : r2_2087;
wire r3_1045;
assign r3_1045 = in[2]? r2_2090 : r2_2089;
wire r3_1046;
assign r3_1046 = in[2]? r2_2092 : r2_2091;
wire r3_1047;
assign r3_1047 = in[2]? r2_2094 : r2_2093;
wire r3_1048;
assign r3_1048 = in[2]? r2_2096 : r2_2095;
wire r3_1049;
assign r3_1049 = in[2]? r2_2098 : r2_2097;
wire r3_1050;
assign r3_1050 = in[2]? r2_2100 : r2_2099;
wire r3_1051;
assign r3_1051 = in[2]? r2_2102 : r2_2101;
wire r3_1052;
assign r3_1052 = in[2]? r2_2104 : r2_2103;
wire r3_1053;
assign r3_1053 = in[2]? r2_2106 : r2_2105;
wire r3_1054;
assign r3_1054 = in[2]? r2_2108 : r2_2107;
wire r3_1055;
assign r3_1055 = in[2]? r2_2110 : r2_2109;
wire r3_1056;
assign r3_1056 = in[2]? r2_2112 : r2_2111;
wire r3_1057;
assign r3_1057 = in[2]? r2_2114 : r2_2113;
wire r3_1058;
assign r3_1058 = in[2]? r2_2116 : r2_2115;
wire r3_1059;
assign r3_1059 = in[2]? r2_2118 : r2_2117;
wire r3_1060;
assign r3_1060 = in[2]? r2_2120 : r2_2119;
wire r3_1061;
assign r3_1061 = in[2]? r2_2122 : r2_2121;
wire r3_1062;
assign r3_1062 = in[2]? r2_2124 : r2_2123;
wire r3_1063;
assign r3_1063 = in[2]? r2_2126 : r2_2125;
wire r3_1064;
assign r3_1064 = in[2]? r2_2128 : r2_2127;
wire r3_1065;
assign r3_1065 = in[2]? r2_2130 : r2_2129;
wire r3_1066;
assign r3_1066 = in[2]? r2_2132 : r2_2131;
wire r3_1067;
assign r3_1067 = in[2]? r2_2134 : r2_2133;
wire r3_1068;
assign r3_1068 = in[2]? r2_2136 : r2_2135;
wire r3_1069;
assign r3_1069 = in[2]? r2_2138 : r2_2137;
wire r3_1070;
assign r3_1070 = in[2]? r2_2140 : r2_2139;
wire r3_1071;
assign r3_1071 = in[2]? r2_2142 : r2_2141;
wire r3_1072;
assign r3_1072 = in[2]? r2_2144 : r2_2143;
wire r3_1073;
assign r3_1073 = in[2]? r2_2146 : r2_2145;
wire r3_1074;
assign r3_1074 = in[2]? r2_2148 : r2_2147;
wire r3_1075;
assign r3_1075 = in[2]? r2_2150 : r2_2149;
wire r3_1076;
assign r3_1076 = in[2]? r2_2152 : r2_2151;
wire r3_1077;
assign r3_1077 = in[2]? r2_2154 : r2_2153;
wire r3_1078;
assign r3_1078 = in[2]? r2_2156 : r2_2155;
wire r3_1079;
assign r3_1079 = in[2]? r2_2158 : r2_2157;
wire r3_1080;
assign r3_1080 = in[2]? r2_2160 : r2_2159;
wire r3_1081;
assign r3_1081 = in[2]? r2_2162 : r2_2161;
wire r3_1082;
assign r3_1082 = in[2]? r2_2164 : r2_2163;
wire r3_1083;
assign r3_1083 = in[2]? r2_2166 : r2_2165;
wire r3_1084;
assign r3_1084 = in[2]? r2_2168 : r2_2167;
wire r3_1085;
assign r3_1085 = in[2]? r2_2170 : r2_2169;
wire r3_1086;
assign r3_1086 = in[2]? r2_2172 : r2_2171;
wire r3_1087;
assign r3_1087 = in[2]? r2_2174 : r2_2173;
wire r3_1088;
assign r3_1088 = in[2]? r2_2176 : r2_2175;
wire r3_1089;
assign r3_1089 = in[2]? r2_2178 : r2_2177;
wire r3_1090;
assign r3_1090 = in[2]? r2_2180 : r2_2179;
wire r3_1091;
assign r3_1091 = in[2]? r2_2182 : r2_2181;
wire r3_1092;
assign r3_1092 = in[2]? r2_2184 : r2_2183;
wire r3_1093;
assign r3_1093 = in[2]? r2_2186 : r2_2185;
wire r3_1094;
assign r3_1094 = in[2]? r2_2188 : r2_2187;
wire r3_1095;
assign r3_1095 = in[2]? r2_2190 : r2_2189;
wire r3_1096;
assign r3_1096 = in[2]? r2_2192 : r2_2191;
wire r3_1097;
assign r3_1097 = in[2]? r2_2194 : r2_2193;
wire r3_1098;
assign r3_1098 = in[2]? r2_2196 : r2_2195;
wire r3_1099;
assign r3_1099 = in[2]? r2_2198 : r2_2197;
wire r3_1100;
assign r3_1100 = in[2]? r2_2200 : r2_2199;
wire r3_1101;
assign r3_1101 = in[2]? r2_2202 : r2_2201;
wire r3_1102;
assign r3_1102 = in[2]? r2_2204 : r2_2203;
wire r3_1103;
assign r3_1103 = in[2]? r2_2206 : r2_2205;
wire r3_1104;
assign r3_1104 = in[2]? r2_2208 : r2_2207;
wire r3_1105;
assign r3_1105 = in[2]? r2_2210 : r2_2209;
wire r3_1106;
assign r3_1106 = in[2]? r2_2212 : r2_2211;
wire r3_1107;
assign r3_1107 = in[2]? r2_2214 : r2_2213;
wire r3_1108;
assign r3_1108 = in[2]? r2_2216 : r2_2215;
wire r3_1109;
assign r3_1109 = in[2]? r2_2218 : r2_2217;
wire r3_1110;
assign r3_1110 = in[2]? r2_2220 : r2_2219;
wire r3_1111;
assign r3_1111 = in[2]? r2_2222 : r2_2221;
wire r3_1112;
assign r3_1112 = in[2]? r2_2224 : r2_2223;
wire r3_1113;
assign r3_1113 = in[2]? r2_2226 : r2_2225;
wire r3_1114;
assign r3_1114 = in[2]? r2_2228 : r2_2227;
wire r3_1115;
assign r3_1115 = in[2]? r2_2230 : r2_2229;
wire r3_1116;
assign r3_1116 = in[2]? r2_2232 : r2_2231;
wire r3_1117;
assign r3_1117 = in[2]? r2_2234 : r2_2233;
wire r3_1118;
assign r3_1118 = in[2]? r2_2236 : r2_2235;
wire r3_1119;
assign r3_1119 = in[2]? r2_2238 : r2_2237;
wire r3_1120;
assign r3_1120 = in[2]? r2_2240 : r2_2239;
wire r3_1121;
assign r3_1121 = in[2]? r2_2242 : r2_2241;
wire r3_1122;
assign r3_1122 = in[2]? r2_2244 : r2_2243;
wire r3_1123;
assign r3_1123 = in[2]? r2_2246 : r2_2245;
wire r3_1124;
assign r3_1124 = in[2]? r2_2248 : r2_2247;
wire r3_1125;
assign r3_1125 = in[2]? r2_2250 : r2_2249;
wire r3_1126;
assign r3_1126 = in[2]? r2_2252 : r2_2251;
wire r3_1127;
assign r3_1127 = in[2]? r2_2254 : r2_2253;
wire r3_1128;
assign r3_1128 = in[2]? r2_2256 : r2_2255;
wire r3_1129;
assign r3_1129 = in[2]? r2_2258 : r2_2257;
wire r3_1130;
assign r3_1130 = in[2]? r2_2260 : r2_2259;
wire r3_1131;
assign r3_1131 = in[2]? r2_2262 : r2_2261;
wire r3_1132;
assign r3_1132 = in[2]? r2_2264 : r2_2263;
wire r3_1133;
assign r3_1133 = in[2]? r2_2266 : r2_2265;
wire r3_1134;
assign r3_1134 = in[2]? r2_2268 : r2_2267;
wire r3_1135;
assign r3_1135 = in[2]? r2_2270 : r2_2269;
wire r3_1136;
assign r3_1136 = in[2]? r2_2272 : r2_2271;
wire r3_1137;
assign r3_1137 = in[2]? r2_2274 : r2_2273;
wire r3_1138;
assign r3_1138 = in[2]? r2_2276 : r2_2275;
wire r3_1139;
assign r3_1139 = in[2]? r2_2278 : r2_2277;
wire r3_1140;
assign r3_1140 = in[2]? r2_2280 : r2_2279;
wire r3_1141;
assign r3_1141 = in[2]? r2_2282 : r2_2281;
wire r3_1142;
assign r3_1142 = in[2]? r2_2284 : r2_2283;
wire r3_1143;
assign r3_1143 = in[2]? r2_2286 : r2_2285;
wire r3_1144;
assign r3_1144 = in[2]? r2_2288 : r2_2287;
wire r3_1145;
assign r3_1145 = in[2]? r2_2290 : r2_2289;
wire r3_1146;
assign r3_1146 = in[2]? r2_2292 : r2_2291;
wire r3_1147;
assign r3_1147 = in[2]? r2_2294 : r2_2293;
wire r3_1148;
assign r3_1148 = in[2]? r2_2296 : r2_2295;
wire r3_1149;
assign r3_1149 = in[2]? r2_2298 : r2_2297;
wire r3_1150;
assign r3_1150 = in[2]? r2_2300 : r2_2299;
wire r3_1151;
assign r3_1151 = in[2]? r2_2302 : r2_2301;
wire r3_1152;
assign r3_1152 = in[2]? r2_2304 : r2_2303;
wire r3_1153;
assign r3_1153 = in[2]? r2_2306 : r2_2305;
wire r3_1154;
assign r3_1154 = in[2]? r2_2308 : r2_2307;
wire r3_1155;
assign r3_1155 = in[2]? r2_2310 : r2_2309;
wire r3_1156;
assign r3_1156 = in[2]? r2_2312 : r2_2311;
wire r3_1157;
assign r3_1157 = in[2]? r2_2314 : r2_2313;
wire r3_1158;
assign r3_1158 = in[2]? r2_2316 : r2_2315;
wire r3_1159;
assign r3_1159 = in[2]? r2_2318 : r2_2317;
wire r3_1160;
assign r3_1160 = in[2]? r2_2320 : r2_2319;
wire r3_1161;
assign r3_1161 = in[2]? r2_2322 : r2_2321;
wire r3_1162;
assign r3_1162 = in[2]? r2_2324 : r2_2323;
wire r3_1163;
assign r3_1163 = in[2]? r2_2326 : r2_2325;
wire r3_1164;
assign r3_1164 = in[2]? r2_2328 : r2_2327;
wire r3_1165;
assign r3_1165 = in[2]? r2_2330 : r2_2329;
wire r3_1166;
assign r3_1166 = in[2]? r2_2332 : r2_2331;
wire r3_1167;
assign r3_1167 = in[2]? r2_2334 : r2_2333;
wire r3_1168;
assign r3_1168 = in[2]? r2_2336 : r2_2335;
wire r3_1169;
assign r3_1169 = in[2]? r2_2338 : r2_2337;
wire r3_1170;
assign r3_1170 = in[2]? r2_2340 : r2_2339;
wire r3_1171;
assign r3_1171 = in[2]? r2_2342 : r2_2341;
wire r3_1172;
assign r3_1172 = in[2]? r2_2344 : r2_2343;
wire r3_1173;
assign r3_1173 = in[2]? r2_2346 : r2_2345;
wire r3_1174;
assign r3_1174 = in[2]? r2_2348 : r2_2347;
wire r3_1175;
assign r3_1175 = in[2]? r2_2350 : r2_2349;
wire r3_1176;
assign r3_1176 = in[2]? r2_2352 : r2_2351;
wire r3_1177;
assign r3_1177 = in[2]? r2_2354 : r2_2353;
wire r3_1178;
assign r3_1178 = in[2]? r2_2356 : r2_2355;
wire r3_1179;
assign r3_1179 = in[2]? r2_2358 : r2_2357;
wire r3_1180;
assign r3_1180 = in[2]? r2_2360 : r2_2359;
wire r3_1181;
assign r3_1181 = in[2]? r2_2362 : r2_2361;
wire r3_1182;
assign r3_1182 = in[2]? r2_2364 : r2_2363;
wire r3_1183;
assign r3_1183 = in[2]? r2_2366 : r2_2365;
wire r3_1184;
assign r3_1184 = in[2]? r2_2368 : r2_2367;
wire r3_1185;
assign r3_1185 = in[2]? r2_2370 : r2_2369;
wire r3_1186;
assign r3_1186 = in[2]? r2_2372 : r2_2371;
wire r3_1187;
assign r3_1187 = in[2]? r2_2374 : r2_2373;
wire r3_1188;
assign r3_1188 = in[2]? r2_2376 : r2_2375;
wire r3_1189;
assign r3_1189 = in[2]? r2_2378 : r2_2377;
wire r3_1190;
assign r3_1190 = in[2]? r2_2380 : r2_2379;
wire r3_1191;
assign r3_1191 = in[2]? r2_2382 : r2_2381;
wire r3_1192;
assign r3_1192 = in[2]? r2_2384 : r2_2383;
wire r3_1193;
assign r3_1193 = in[2]? r2_2386 : r2_2385;
wire r3_1194;
assign r3_1194 = in[2]? r2_2388 : r2_2387;
wire r3_1195;
assign r3_1195 = in[2]? r2_2390 : r2_2389;
wire r3_1196;
assign r3_1196 = in[2]? r2_2392 : r2_2391;
wire r3_1197;
assign r3_1197 = in[2]? r2_2394 : r2_2393;
wire r3_1198;
assign r3_1198 = in[2]? r2_2396 : r2_2395;
wire r3_1199;
assign r3_1199 = in[2]? r2_2398 : r2_2397;
wire r3_1200;
assign r3_1200 = in[2]? r2_2400 : r2_2399;
wire r3_1201;
assign r3_1201 = in[2]? r2_2402 : r2_2401;
wire r3_1202;
assign r3_1202 = in[2]? r2_2404 : r2_2403;
wire r3_1203;
assign r3_1203 = in[2]? r2_2406 : r2_2405;
wire r3_1204;
assign r3_1204 = in[2]? r2_2408 : r2_2407;
wire r3_1205;
assign r3_1205 = in[2]? r2_2410 : r2_2409;
wire r3_1206;
assign r3_1206 = in[2]? r2_2412 : r2_2411;
wire r3_1207;
assign r3_1207 = in[2]? r2_2414 : r2_2413;
wire r3_1208;
assign r3_1208 = in[2]? r2_2416 : r2_2415;
wire r3_1209;
assign r3_1209 = in[2]? r2_2418 : r2_2417;
wire r3_1210;
assign r3_1210 = in[2]? r2_2420 : r2_2419;
wire r3_1211;
assign r3_1211 = in[2]? r2_2422 : r2_2421;
wire r3_1212;
assign r3_1212 = in[2]? r2_2424 : r2_2423;
wire r3_1213;
assign r3_1213 = in[2]? r2_2426 : r2_2425;
wire r3_1214;
assign r3_1214 = in[2]? r2_2428 : r2_2427;
wire r3_1215;
assign r3_1215 = in[2]? r2_2430 : r2_2429;
wire r3_1216;
assign r3_1216 = in[2]? r2_2432 : r2_2431;
wire r3_1217;
assign r3_1217 = in[2]? r2_2434 : r2_2433;
wire r3_1218;
assign r3_1218 = in[2]? r2_2436 : r2_2435;
wire r3_1219;
assign r3_1219 = in[2]? r2_2438 : r2_2437;
wire r3_1220;
assign r3_1220 = in[2]? r2_2440 : r2_2439;
wire r3_1221;
assign r3_1221 = in[2]? r2_2442 : r2_2441;
wire r3_1222;
assign r3_1222 = in[2]? r2_2444 : r2_2443;
wire r3_1223;
assign r3_1223 = in[2]? r2_2446 : r2_2445;
wire r3_1224;
assign r3_1224 = in[2]? r2_2448 : r2_2447;
wire r3_1225;
assign r3_1225 = in[2]? r2_2450 : r2_2449;
wire r3_1226;
assign r3_1226 = in[2]? r2_2452 : r2_2451;
wire r3_1227;
assign r3_1227 = in[2]? r2_2454 : r2_2453;
wire r3_1228;
assign r3_1228 = in[2]? r2_2456 : r2_2455;
wire r3_1229;
assign r3_1229 = in[2]? r2_2458 : r2_2457;
wire r3_1230;
assign r3_1230 = in[2]? r2_2460 : r2_2459;
wire r3_1231;
assign r3_1231 = in[2]? r2_2462 : r2_2461;
wire r3_1232;
assign r3_1232 = in[2]? r2_2464 : r2_2463;
wire r3_1233;
assign r3_1233 = in[2]? r2_2466 : r2_2465;
wire r3_1234;
assign r3_1234 = in[2]? r2_2468 : r2_2467;
wire r3_1235;
assign r3_1235 = in[2]? r2_2470 : r2_2469;
wire r3_1236;
assign r3_1236 = in[2]? r2_2472 : r2_2471;
wire r3_1237;
assign r3_1237 = in[2]? r2_2474 : r2_2473;
wire r3_1238;
assign r3_1238 = in[2]? r2_2476 : r2_2475;
wire r3_1239;
assign r3_1239 = in[2]? r2_2478 : r2_2477;
wire r3_1240;
assign r3_1240 = in[2]? r2_2480 : r2_2479;
wire r3_1241;
assign r3_1241 = in[2]? r2_2482 : r2_2481;
wire r3_1242;
assign r3_1242 = in[2]? r2_2484 : r2_2483;
wire r3_1243;
assign r3_1243 = in[2]? r2_2486 : r2_2485;
wire r3_1244;
assign r3_1244 = in[2]? r2_2488 : r2_2487;
wire r3_1245;
assign r3_1245 = in[2]? r2_2490 : r2_2489;
wire r3_1246;
assign r3_1246 = in[2]? r2_2492 : r2_2491;
wire r3_1247;
assign r3_1247 = in[2]? r2_2494 : r2_2493;
wire r3_1248;
assign r3_1248 = in[2]? r2_2496 : r2_2495;
wire r3_1249;
assign r3_1249 = in[2]? r2_2498 : r2_2497;
wire r3_1250;
assign r3_1250 = in[2]? r2_2500 : r2_2499;
wire r3_1251;
assign r3_1251 = in[2]? r2_2502 : r2_2501;
wire r3_1252;
assign r3_1252 = in[2]? r2_2504 : r2_2503;
wire r3_1253;
assign r3_1253 = in[2]? r2_2506 : r2_2505;
wire r3_1254;
assign r3_1254 = in[2]? r2_2508 : r2_2507;
wire r3_1255;
assign r3_1255 = in[2]? r2_2510 : r2_2509;
wire r3_1256;
assign r3_1256 = in[2]? r2_2512 : r2_2511;
wire r3_1257;
assign r3_1257 = in[2]? r2_2514 : r2_2513;
wire r3_1258;
assign r3_1258 = in[2]? r2_2516 : r2_2515;
wire r3_1259;
assign r3_1259 = in[2]? r2_2518 : r2_2517;
wire r3_1260;
assign r3_1260 = in[2]? r2_2520 : r2_2519;
wire r3_1261;
assign r3_1261 = in[2]? r2_2522 : r2_2521;
wire r3_1262;
assign r3_1262 = in[2]? r2_2524 : r2_2523;
wire r3_1263;
assign r3_1263 = in[2]? r2_2526 : r2_2525;
wire r3_1264;
assign r3_1264 = in[2]? r2_2528 : r2_2527;
wire r3_1265;
assign r3_1265 = in[2]? r2_2530 : r2_2529;
wire r3_1266;
assign r3_1266 = in[2]? r2_2532 : r2_2531;
wire r3_1267;
assign r3_1267 = in[2]? r2_2534 : r2_2533;
wire r3_1268;
assign r3_1268 = in[2]? r2_2536 : r2_2535;
wire r3_1269;
assign r3_1269 = in[2]? r2_2538 : r2_2537;
wire r3_1270;
assign r3_1270 = in[2]? r2_2540 : r2_2539;
wire r3_1271;
assign r3_1271 = in[2]? r2_2542 : r2_2541;
wire r3_1272;
assign r3_1272 = in[2]? r2_2544 : r2_2543;
wire r3_1273;
assign r3_1273 = in[2]? r2_2546 : r2_2545;
wire r3_1274;
assign r3_1274 = in[2]? r2_2548 : r2_2547;
wire r3_1275;
assign r3_1275 = in[2]? r2_2550 : r2_2549;
wire r3_1276;
assign r3_1276 = in[2]? r2_2552 : r2_2551;
wire r3_1277;
assign r3_1277 = in[2]? r2_2554 : r2_2553;
wire r3_1278;
assign r3_1278 = in[2]? r2_2556 : r2_2555;
wire r3_1279;
assign r3_1279 = in[2]? r2_2558 : r2_2557;
wire r3_1280;
assign r3_1280 = in[2]? r2_2560 : r2_2559;
wire r3_1281;
assign r3_1281 = in[2]? r2_2562 : r2_2561;
wire r3_1282;
assign r3_1282 = in[2]? r2_2564 : r2_2563;
wire r3_1283;
assign r3_1283 = in[2]? r2_2566 : r2_2565;
wire r3_1284;
assign r3_1284 = in[2]? r2_2568 : r2_2567;
wire r3_1285;
assign r3_1285 = in[2]? r2_2570 : r2_2569;
wire r3_1286;
assign r3_1286 = in[2]? r2_2572 : r2_2571;
wire r3_1287;
assign r3_1287 = in[2]? r2_2574 : r2_2573;
wire r3_1288;
assign r3_1288 = in[2]? r2_2576 : r2_2575;
wire r3_1289;
assign r3_1289 = in[2]? r2_2578 : r2_2577;
wire r3_1290;
assign r3_1290 = in[2]? r2_2580 : r2_2579;
wire r3_1291;
assign r3_1291 = in[2]? r2_2582 : r2_2581;
wire r3_1292;
assign r3_1292 = in[2]? r2_2584 : r2_2583;
wire r3_1293;
assign r3_1293 = in[2]? r2_2586 : r2_2585;
wire r3_1294;
assign r3_1294 = in[2]? r2_2588 : r2_2587;
wire r3_1295;
assign r3_1295 = in[2]? r2_2590 : r2_2589;
wire r3_1296;
assign r3_1296 = in[2]? r2_2592 : r2_2591;
wire r3_1297;
assign r3_1297 = in[2]? r2_2594 : r2_2593;
wire r3_1298;
assign r3_1298 = in[2]? r2_2596 : r2_2595;
wire r3_1299;
assign r3_1299 = in[2]? r2_2598 : r2_2597;
wire r3_1300;
assign r3_1300 = in[2]? r2_2600 : r2_2599;
wire r3_1301;
assign r3_1301 = in[2]? r2_2602 : r2_2601;
wire r3_1302;
assign r3_1302 = in[2]? r2_2604 : r2_2603;
wire r3_1303;
assign r3_1303 = in[2]? r2_2606 : r2_2605;
wire r3_1304;
assign r3_1304 = in[2]? r2_2608 : r2_2607;
wire r3_1305;
assign r3_1305 = in[2]? r2_2610 : r2_2609;
wire r3_1306;
assign r3_1306 = in[2]? r2_2612 : r2_2611;
wire r3_1307;
assign r3_1307 = in[2]? r2_2614 : r2_2613;
wire r3_1308;
assign r3_1308 = in[2]? r2_2616 : r2_2615;
wire r3_1309;
assign r3_1309 = in[2]? r2_2618 : r2_2617;
wire r3_1310;
assign r3_1310 = in[2]? r2_2620 : r2_2619;
wire r3_1311;
assign r3_1311 = in[2]? r2_2622 : r2_2621;
wire r3_1312;
assign r3_1312 = in[2]? r2_2624 : r2_2623;
wire r3_1313;
assign r3_1313 = in[2]? r2_2626 : r2_2625;
wire r3_1314;
assign r3_1314 = in[2]? r2_2628 : r2_2627;
wire r3_1315;
assign r3_1315 = in[2]? r2_2630 : r2_2629;
wire r3_1316;
assign r3_1316 = in[2]? r2_2632 : r2_2631;
wire r3_1317;
assign r3_1317 = in[2]? r2_2634 : r2_2633;
wire r3_1318;
assign r3_1318 = in[2]? r2_2636 : r2_2635;
wire r3_1319;
assign r3_1319 = in[2]? r2_2638 : r2_2637;
wire r3_1320;
assign r3_1320 = in[2]? r2_2640 : r2_2639;
wire r3_1321;
assign r3_1321 = in[2]? r2_2642 : r2_2641;
wire r3_1322;
assign r3_1322 = in[2]? r2_2644 : r2_2643;
wire r3_1323;
assign r3_1323 = in[2]? r2_2646 : r2_2645;
wire r3_1324;
assign r3_1324 = in[2]? r2_2648 : r2_2647;
wire r3_1325;
assign r3_1325 = in[2]? r2_2650 : r2_2649;
wire r3_1326;
assign r3_1326 = in[2]? r2_2652 : r2_2651;
wire r3_1327;
assign r3_1327 = in[2]? r2_2654 : r2_2653;
wire r3_1328;
assign r3_1328 = in[2]? r2_2656 : r2_2655;
wire r3_1329;
assign r3_1329 = in[2]? r2_2658 : r2_2657;
wire r3_1330;
assign r3_1330 = in[2]? r2_2660 : r2_2659;
wire r3_1331;
assign r3_1331 = in[2]? r2_2662 : r2_2661;
wire r3_1332;
assign r3_1332 = in[2]? r2_2664 : r2_2663;
wire r3_1333;
assign r3_1333 = in[2]? r2_2666 : r2_2665;
wire r3_1334;
assign r3_1334 = in[2]? r2_2668 : r2_2667;
wire r3_1335;
assign r3_1335 = in[2]? r2_2670 : r2_2669;
wire r3_1336;
assign r3_1336 = in[2]? r2_2672 : r2_2671;
wire r3_1337;
assign r3_1337 = in[2]? r2_2674 : r2_2673;
wire r3_1338;
assign r3_1338 = in[2]? r2_2676 : r2_2675;
wire r3_1339;
assign r3_1339 = in[2]? r2_2678 : r2_2677;
wire r3_1340;
assign r3_1340 = in[2]? r2_2680 : r2_2679;
wire r3_1341;
assign r3_1341 = in[2]? r2_2682 : r2_2681;
wire r3_1342;
assign r3_1342 = in[2]? r2_2684 : r2_2683;
wire r3_1343;
assign r3_1343 = in[2]? r2_2686 : r2_2685;
wire r3_1344;
assign r3_1344 = in[2]? r2_2688 : r2_2687;
wire r3_1345;
assign r3_1345 = in[2]? r2_2690 : r2_2689;
wire r3_1346;
assign r3_1346 = in[2]? r2_2692 : r2_2691;
wire r3_1347;
assign r3_1347 = in[2]? r2_2694 : r2_2693;
wire r3_1348;
assign r3_1348 = in[2]? r2_2696 : r2_2695;
wire r3_1349;
assign r3_1349 = in[2]? r2_2698 : r2_2697;
wire r3_1350;
assign r3_1350 = in[2]? r2_2700 : r2_2699;
wire r3_1351;
assign r3_1351 = in[2]? r2_2702 : r2_2701;
wire r3_1352;
assign r3_1352 = in[2]? r2_2704 : r2_2703;
wire r3_1353;
assign r3_1353 = in[2]? r2_2706 : r2_2705;
wire r3_1354;
assign r3_1354 = in[2]? r2_2708 : r2_2707;
wire r3_1355;
assign r3_1355 = in[2]? r2_2710 : r2_2709;
wire r3_1356;
assign r3_1356 = in[2]? r2_2712 : r2_2711;
wire r3_1357;
assign r3_1357 = in[2]? r2_2714 : r2_2713;
wire r3_1358;
assign r3_1358 = in[2]? r2_2716 : r2_2715;
wire r3_1359;
assign r3_1359 = in[2]? r2_2718 : r2_2717;
wire r3_1360;
assign r3_1360 = in[2]? r2_2720 : r2_2719;
wire r3_1361;
assign r3_1361 = in[2]? r2_2722 : r2_2721;
wire r3_1362;
assign r3_1362 = in[2]? r2_2724 : r2_2723;
wire r3_1363;
assign r3_1363 = in[2]? r2_2726 : r2_2725;
wire r3_1364;
assign r3_1364 = in[2]? r2_2728 : r2_2727;
wire r3_1365;
assign r3_1365 = in[2]? r2_2730 : r2_2729;
wire r3_1366;
assign r3_1366 = in[2]? r2_2732 : r2_2731;
wire r3_1367;
assign r3_1367 = in[2]? r2_2734 : r2_2733;
wire r3_1368;
assign r3_1368 = in[2]? r2_2736 : r2_2735;
wire r3_1369;
assign r3_1369 = in[2]? r2_2738 : r2_2737;
wire r3_1370;
assign r3_1370 = in[2]? r2_2740 : r2_2739;
wire r3_1371;
assign r3_1371 = in[2]? r2_2742 : r2_2741;
wire r3_1372;
assign r3_1372 = in[2]? r2_2744 : r2_2743;
wire r3_1373;
assign r3_1373 = in[2]? r2_2746 : r2_2745;
wire r3_1374;
assign r3_1374 = in[2]? r2_2748 : r2_2747;
wire r3_1375;
assign r3_1375 = in[2]? r2_2750 : r2_2749;
wire r3_1376;
assign r3_1376 = in[2]? r2_2752 : r2_2751;
wire r3_1377;
assign r3_1377 = in[2]? r2_2754 : r2_2753;
wire r3_1378;
assign r3_1378 = in[2]? r2_2756 : r2_2755;
wire r3_1379;
assign r3_1379 = in[2]? r2_2758 : r2_2757;
wire r3_1380;
assign r3_1380 = in[2]? r2_2760 : r2_2759;
wire r3_1381;
assign r3_1381 = in[2]? r2_2762 : r2_2761;
wire r3_1382;
assign r3_1382 = in[2]? r2_2764 : r2_2763;
wire r3_1383;
assign r3_1383 = in[2]? r2_2766 : r2_2765;
wire r3_1384;
assign r3_1384 = in[2]? r2_2768 : r2_2767;
wire r3_1385;
assign r3_1385 = in[2]? r2_2770 : r2_2769;
wire r3_1386;
assign r3_1386 = in[2]? r2_2772 : r2_2771;
wire r3_1387;
assign r3_1387 = in[2]? r2_2774 : r2_2773;
wire r3_1388;
assign r3_1388 = in[2]? r2_2776 : r2_2775;
wire r3_1389;
assign r3_1389 = in[2]? r2_2778 : r2_2777;
wire r3_1390;
assign r3_1390 = in[2]? r2_2780 : r2_2779;
wire r3_1391;
assign r3_1391 = in[2]? r2_2782 : r2_2781;
wire r3_1392;
assign r3_1392 = in[2]? r2_2784 : r2_2783;
wire r3_1393;
assign r3_1393 = in[2]? r2_2786 : r2_2785;
wire r3_1394;
assign r3_1394 = in[2]? r2_2788 : r2_2787;
wire r3_1395;
assign r3_1395 = in[2]? r2_2790 : r2_2789;
wire r3_1396;
assign r3_1396 = in[2]? r2_2792 : r2_2791;
wire r3_1397;
assign r3_1397 = in[2]? r2_2794 : r2_2793;
wire r3_1398;
assign r3_1398 = in[2]? r2_2796 : r2_2795;
wire r3_1399;
assign r3_1399 = in[2]? r2_2798 : r2_2797;
wire r3_1400;
assign r3_1400 = in[2]? r2_2800 : r2_2799;
wire r3_1401;
assign r3_1401 = in[2]? r2_2802 : r2_2801;
wire r3_1402;
assign r3_1402 = in[2]? r2_2804 : r2_2803;
wire r3_1403;
assign r3_1403 = in[2]? r2_2806 : r2_2805;
wire r3_1404;
assign r3_1404 = in[2]? r2_2808 : r2_2807;
wire r3_1405;
assign r3_1405 = in[2]? r2_2810 : r2_2809;
wire r3_1406;
assign r3_1406 = in[2]? r2_2812 : r2_2811;
wire r3_1407;
assign r3_1407 = in[2]? r2_2814 : r2_2813;
wire r3_1408;
assign r3_1408 = in[2]? r2_2816 : r2_2815;
wire r3_1409;
assign r3_1409 = in[2]? r2_2818 : r2_2817;
wire r3_1410;
assign r3_1410 = in[2]? r2_2820 : r2_2819;
wire r3_1411;
assign r3_1411 = in[2]? r2_2822 : r2_2821;
wire r3_1412;
assign r3_1412 = in[2]? r2_2824 : r2_2823;
wire r3_1413;
assign r3_1413 = in[2]? r2_2826 : r2_2825;
wire r3_1414;
assign r3_1414 = in[2]? r2_2828 : r2_2827;
wire r3_1415;
assign r3_1415 = in[2]? r2_2830 : r2_2829;
wire r3_1416;
assign r3_1416 = in[2]? r2_2832 : r2_2831;
wire r3_1417;
assign r3_1417 = in[2]? r2_2834 : r2_2833;
wire r3_1418;
assign r3_1418 = in[2]? r2_2836 : r2_2835;
wire r3_1419;
assign r3_1419 = in[2]? r2_2838 : r2_2837;
wire r3_1420;
assign r3_1420 = in[2]? r2_2840 : r2_2839;
wire r3_1421;
assign r3_1421 = in[2]? r2_2842 : r2_2841;
wire r3_1422;
assign r3_1422 = in[2]? r2_2844 : r2_2843;
wire r3_1423;
assign r3_1423 = in[2]? r2_2846 : r2_2845;
wire r3_1424;
assign r3_1424 = in[2]? r2_2848 : r2_2847;
wire r3_1425;
assign r3_1425 = in[2]? r2_2850 : r2_2849;
wire r3_1426;
assign r3_1426 = in[2]? r2_2852 : r2_2851;
wire r3_1427;
assign r3_1427 = in[2]? r2_2854 : r2_2853;
wire r3_1428;
assign r3_1428 = in[2]? r2_2856 : r2_2855;
wire r3_1429;
assign r3_1429 = in[2]? r2_2858 : r2_2857;
wire r3_1430;
assign r3_1430 = in[2]? r2_2860 : r2_2859;
wire r3_1431;
assign r3_1431 = in[2]? r2_2862 : r2_2861;
wire r3_1432;
assign r3_1432 = in[2]? r2_2864 : r2_2863;
wire r3_1433;
assign r3_1433 = in[2]? r2_2866 : r2_2865;
wire r3_1434;
assign r3_1434 = in[2]? r2_2868 : r2_2867;
wire r3_1435;
assign r3_1435 = in[2]? r2_2870 : r2_2869;
wire r3_1436;
assign r3_1436 = in[2]? r2_2872 : r2_2871;
wire r3_1437;
assign r3_1437 = in[2]? r2_2874 : r2_2873;
wire r3_1438;
assign r3_1438 = in[2]? r2_2876 : r2_2875;
wire r3_1439;
assign r3_1439 = in[2]? r2_2878 : r2_2877;
wire r3_1440;
assign r3_1440 = in[2]? r2_2880 : r2_2879;
wire r3_1441;
assign r3_1441 = in[2]? r2_2882 : r2_2881;
wire r3_1442;
assign r3_1442 = in[2]? r2_2884 : r2_2883;
wire r3_1443;
assign r3_1443 = in[2]? r2_2886 : r2_2885;
wire r3_1444;
assign r3_1444 = in[2]? r2_2888 : r2_2887;
wire r3_1445;
assign r3_1445 = in[2]? r2_2890 : r2_2889;
wire r3_1446;
assign r3_1446 = in[2]? r2_2892 : r2_2891;
wire r3_1447;
assign r3_1447 = in[2]? r2_2894 : r2_2893;
wire r3_1448;
assign r3_1448 = in[2]? r2_2896 : r2_2895;
wire r3_1449;
assign r3_1449 = in[2]? r2_2898 : r2_2897;
wire r3_1450;
assign r3_1450 = in[2]? r2_2900 : r2_2899;
wire r3_1451;
assign r3_1451 = in[2]? r2_2902 : r2_2901;
wire r3_1452;
assign r3_1452 = in[2]? r2_2904 : r2_2903;
wire r3_1453;
assign r3_1453 = in[2]? r2_2906 : r2_2905;
wire r3_1454;
assign r3_1454 = in[2]? r2_2908 : r2_2907;
wire r3_1455;
assign r3_1455 = in[2]? r2_2910 : r2_2909;
wire r3_1456;
assign r3_1456 = in[2]? r2_2912 : r2_2911;
wire r3_1457;
assign r3_1457 = in[2]? r2_2914 : r2_2913;
wire r3_1458;
assign r3_1458 = in[2]? r2_2916 : r2_2915;
wire r3_1459;
assign r3_1459 = in[2]? r2_2918 : r2_2917;
wire r3_1460;
assign r3_1460 = in[2]? r2_2920 : r2_2919;
wire r3_1461;
assign r3_1461 = in[2]? r2_2922 : r2_2921;
wire r3_1462;
assign r3_1462 = in[2]? r2_2924 : r2_2923;
wire r3_1463;
assign r3_1463 = in[2]? r2_2926 : r2_2925;
wire r3_1464;
assign r3_1464 = in[2]? r2_2928 : r2_2927;
wire r3_1465;
assign r3_1465 = in[2]? r2_2930 : r2_2929;
wire r3_1466;
assign r3_1466 = in[2]? r2_2932 : r2_2931;
wire r3_1467;
assign r3_1467 = in[2]? r2_2934 : r2_2933;
wire r3_1468;
assign r3_1468 = in[2]? r2_2936 : r2_2935;
wire r3_1469;
assign r3_1469 = in[2]? r2_2938 : r2_2937;
wire r3_1470;
assign r3_1470 = in[2]? r2_2940 : r2_2939;
wire r3_1471;
assign r3_1471 = in[2]? r2_2942 : r2_2941;
wire r3_1472;
assign r3_1472 = in[2]? r2_2944 : r2_2943;
wire r3_1473;
assign r3_1473 = in[2]? r2_2946 : r2_2945;
wire r3_1474;
assign r3_1474 = in[2]? r2_2948 : r2_2947;
wire r3_1475;
assign r3_1475 = in[2]? r2_2950 : r2_2949;
wire r3_1476;
assign r3_1476 = in[2]? r2_2952 : r2_2951;
wire r3_1477;
assign r3_1477 = in[2]? r2_2954 : r2_2953;
wire r3_1478;
assign r3_1478 = in[2]? r2_2956 : r2_2955;
wire r3_1479;
assign r3_1479 = in[2]? r2_2958 : r2_2957;
wire r3_1480;
assign r3_1480 = in[2]? r2_2960 : r2_2959;
wire r3_1481;
assign r3_1481 = in[2]? r2_2962 : r2_2961;
wire r3_1482;
assign r3_1482 = in[2]? r2_2964 : r2_2963;
wire r3_1483;
assign r3_1483 = in[2]? r2_2966 : r2_2965;
wire r3_1484;
assign r3_1484 = in[2]? r2_2968 : r2_2967;
wire r3_1485;
assign r3_1485 = in[2]? r2_2970 : r2_2969;
wire r3_1486;
assign r3_1486 = in[2]? r2_2972 : r2_2971;
wire r3_1487;
assign r3_1487 = in[2]? r2_2974 : r2_2973;
wire r3_1488;
assign r3_1488 = in[2]? r2_2976 : r2_2975;
wire r3_1489;
assign r3_1489 = in[2]? r2_2978 : r2_2977;
wire r3_1490;
assign r3_1490 = in[2]? r2_2980 : r2_2979;
wire r3_1491;
assign r3_1491 = in[2]? r2_2982 : r2_2981;
wire r3_1492;
assign r3_1492 = in[2]? r2_2984 : r2_2983;
wire r3_1493;
assign r3_1493 = in[2]? r2_2986 : r2_2985;
wire r3_1494;
assign r3_1494 = in[2]? r2_2988 : r2_2987;
wire r3_1495;
assign r3_1495 = in[2]? r2_2990 : r2_2989;
wire r3_1496;
assign r3_1496 = in[2]? r2_2992 : r2_2991;
wire r3_1497;
assign r3_1497 = in[2]? r2_2994 : r2_2993;
wire r3_1498;
assign r3_1498 = in[2]? r2_2996 : r2_2995;
wire r3_1499;
assign r3_1499 = in[2]? r2_2998 : r2_2997;
wire r3_1500;
assign r3_1500 = in[2]? r2_3000 : r2_2999;
wire r3_1501;
assign r3_1501 = in[2]? r2_3002 : r2_3001;
wire r3_1502;
assign r3_1502 = in[2]? r2_3004 : r2_3003;
wire r3_1503;
assign r3_1503 = in[2]? r2_3006 : r2_3005;
wire r3_1504;
assign r3_1504 = in[2]? r2_3008 : r2_3007;
wire r3_1505;
assign r3_1505 = in[2]? r2_3010 : r2_3009;
wire r3_1506;
assign r3_1506 = in[2]? r2_3012 : r2_3011;
wire r3_1507;
assign r3_1507 = in[2]? r2_3014 : r2_3013;
wire r3_1508;
assign r3_1508 = in[2]? r2_3016 : r2_3015;
wire r3_1509;
assign r3_1509 = in[2]? r2_3018 : r2_3017;
wire r3_1510;
assign r3_1510 = in[2]? r2_3020 : r2_3019;
wire r3_1511;
assign r3_1511 = in[2]? r2_3022 : r2_3021;
wire r3_1512;
assign r3_1512 = in[2]? r2_3024 : r2_3023;
wire r3_1513;
assign r3_1513 = in[2]? r2_3026 : r2_3025;
wire r3_1514;
assign r3_1514 = in[2]? r2_3028 : r2_3027;
wire r3_1515;
assign r3_1515 = in[2]? r2_3030 : r2_3029;
wire r3_1516;
assign r3_1516 = in[2]? r2_3032 : r2_3031;
wire r3_1517;
assign r3_1517 = in[2]? r2_3034 : r2_3033;
wire r3_1518;
assign r3_1518 = in[2]? r2_3036 : r2_3035;
wire r3_1519;
assign r3_1519 = in[2]? r2_3038 : r2_3037;
wire r3_1520;
assign r3_1520 = in[2]? r2_3040 : r2_3039;
wire r3_1521;
assign r3_1521 = in[2]? r2_3042 : r2_3041;
wire r3_1522;
assign r3_1522 = in[2]? r2_3044 : r2_3043;
wire r3_1523;
assign r3_1523 = in[2]? r2_3046 : r2_3045;
wire r3_1524;
assign r3_1524 = in[2]? r2_3048 : r2_3047;
wire r3_1525;
assign r3_1525 = in[2]? r2_3050 : r2_3049;
wire r3_1526;
assign r3_1526 = in[2]? r2_3052 : r2_3051;
wire r3_1527;
assign r3_1527 = in[2]? r2_3054 : r2_3053;
wire r3_1528;
assign r3_1528 = in[2]? r2_3056 : r2_3055;
wire r3_1529;
assign r3_1529 = in[2]? r2_3058 : r2_3057;
wire r3_1530;
assign r3_1530 = in[2]? r2_3060 : r2_3059;
wire r3_1531;
assign r3_1531 = in[2]? r2_3062 : r2_3061;
wire r3_1532;
assign r3_1532 = in[2]? r2_3064 : r2_3063;
wire r3_1533;
assign r3_1533 = in[2]? r2_3066 : r2_3065;
wire r3_1534;
assign r3_1534 = in[2]? r2_3068 : r2_3067;
wire r3_1535;
assign r3_1535 = in[2]? r2_3070 : r2_3069;
wire r3_1536;
assign r3_1536 = in[2]? r2_3072 : r2_3071;
wire r3_1537;
assign r3_1537 = in[2]? r2_3074 : r2_3073;
wire r3_1538;
assign r3_1538 = in[2]? r2_3076 : r2_3075;
wire r3_1539;
assign r3_1539 = in[2]? r2_3078 : r2_3077;
wire r3_1540;
assign r3_1540 = in[2]? r2_3080 : r2_3079;
wire r3_1541;
assign r3_1541 = in[2]? r2_3082 : r2_3081;
wire r3_1542;
assign r3_1542 = in[2]? r2_3084 : r2_3083;
wire r3_1543;
assign r3_1543 = in[2]? r2_3086 : r2_3085;
wire r3_1544;
assign r3_1544 = in[2]? r2_3088 : r2_3087;
wire r3_1545;
assign r3_1545 = in[2]? r2_3090 : r2_3089;
wire r3_1546;
assign r3_1546 = in[2]? r2_3092 : r2_3091;
wire r3_1547;
assign r3_1547 = in[2]? r2_3094 : r2_3093;
wire r3_1548;
assign r3_1548 = in[2]? r2_3096 : r2_3095;
wire r3_1549;
assign r3_1549 = in[2]? r2_3098 : r2_3097;
wire r3_1550;
assign r3_1550 = in[2]? r2_3100 : r2_3099;
wire r3_1551;
assign r3_1551 = in[2]? r2_3102 : r2_3101;
wire r3_1552;
assign r3_1552 = in[2]? r2_3104 : r2_3103;
wire r3_1553;
assign r3_1553 = in[2]? r2_3106 : r2_3105;
wire r3_1554;
assign r3_1554 = in[2]? r2_3108 : r2_3107;
wire r3_1555;
assign r3_1555 = in[2]? r2_3110 : r2_3109;
wire r3_1556;
assign r3_1556 = in[2]? r2_3112 : r2_3111;
wire r3_1557;
assign r3_1557 = in[2]? r2_3114 : r2_3113;
wire r3_1558;
assign r3_1558 = in[2]? r2_3116 : r2_3115;
wire r3_1559;
assign r3_1559 = in[2]? r2_3118 : r2_3117;
wire r3_1560;
assign r3_1560 = in[2]? r2_3120 : r2_3119;
wire r3_1561;
assign r3_1561 = in[2]? r2_3122 : r2_3121;
wire r3_1562;
assign r3_1562 = in[2]? r2_3124 : r2_3123;
wire r3_1563;
assign r3_1563 = in[2]? r2_3126 : r2_3125;
wire r3_1564;
assign r3_1564 = in[2]? r2_3128 : r2_3127;
wire r3_1565;
assign r3_1565 = in[2]? r2_3130 : r2_3129;
wire r3_1566;
assign r3_1566 = in[2]? r2_3132 : r2_3131;
wire r3_1567;
assign r3_1567 = in[2]? r2_3134 : r2_3133;
wire r3_1568;
assign r3_1568 = in[2]? r2_3136 : r2_3135;
wire r3_1569;
assign r3_1569 = in[2]? r2_3138 : r2_3137;
wire r3_1570;
assign r3_1570 = in[2]? r2_3140 : r2_3139;
wire r3_1571;
assign r3_1571 = in[2]? r2_3142 : r2_3141;
wire r3_1572;
assign r3_1572 = in[2]? r2_3144 : r2_3143;
wire r3_1573;
assign r3_1573 = in[2]? r2_3146 : r2_3145;
wire r3_1574;
assign r3_1574 = in[2]? r2_3148 : r2_3147;
wire r3_1575;
assign r3_1575 = in[2]? r2_3150 : r2_3149;
wire r3_1576;
assign r3_1576 = in[2]? r2_3152 : r2_3151;
wire r3_1577;
assign r3_1577 = in[2]? r2_3154 : r2_3153;
wire r3_1578;
assign r3_1578 = in[2]? r2_3156 : r2_3155;
wire r3_1579;
assign r3_1579 = in[2]? r2_3158 : r2_3157;
wire r3_1580;
assign r3_1580 = in[2]? r2_3160 : r2_3159;
wire r3_1581;
assign r3_1581 = in[2]? r2_3162 : r2_3161;
wire r3_1582;
assign r3_1582 = in[2]? r2_3164 : r2_3163;
wire r3_1583;
assign r3_1583 = in[2]? r2_3166 : r2_3165;
wire r3_1584;
assign r3_1584 = in[2]? r2_3168 : r2_3167;
wire r3_1585;
assign r3_1585 = in[2]? r2_3170 : r2_3169;
wire r3_1586;
assign r3_1586 = in[2]? r2_3172 : r2_3171;
wire r3_1587;
assign r3_1587 = in[2]? r2_3174 : r2_3173;
wire r3_1588;
assign r3_1588 = in[2]? r2_3176 : r2_3175;
wire r3_1589;
assign r3_1589 = in[2]? r2_3178 : r2_3177;
wire r3_1590;
assign r3_1590 = in[2]? r2_3180 : r2_3179;
wire r3_1591;
assign r3_1591 = in[2]? r2_3182 : r2_3181;
wire r3_1592;
assign r3_1592 = in[2]? r2_3184 : r2_3183;
wire r3_1593;
assign r3_1593 = in[2]? r2_3186 : r2_3185;
wire r3_1594;
assign r3_1594 = in[2]? r2_3188 : r2_3187;
wire r3_1595;
assign r3_1595 = in[2]? r2_3190 : r2_3189;
wire r3_1596;
assign r3_1596 = in[2]? r2_3192 : r2_3191;
wire r3_1597;
assign r3_1597 = in[2]? r2_3194 : r2_3193;
wire r3_1598;
assign r3_1598 = in[2]? r2_3196 : r2_3195;
wire r3_1599;
assign r3_1599 = in[2]? r2_3198 : r2_3197;
wire r3_1600;
assign r3_1600 = in[2]? r2_3200 : r2_3199;
wire r3_1601;
assign r3_1601 = in[2]? r2_3202 : r2_3201;
wire r3_1602;
assign r3_1602 = in[2]? r2_3204 : r2_3203;
wire r3_1603;
assign r3_1603 = in[2]? r2_3206 : r2_3205;
wire r3_1604;
assign r3_1604 = in[2]? r2_3208 : r2_3207;
wire r3_1605;
assign r3_1605 = in[2]? r2_3210 : r2_3209;
wire r3_1606;
assign r3_1606 = in[2]? r2_3212 : r2_3211;
wire r3_1607;
assign r3_1607 = in[2]? r2_3214 : r2_3213;
wire r3_1608;
assign r3_1608 = in[2]? r2_3216 : r2_3215;
wire r3_1609;
assign r3_1609 = in[2]? r2_3218 : r2_3217;
wire r3_1610;
assign r3_1610 = in[2]? r2_3220 : r2_3219;
wire r3_1611;
assign r3_1611 = in[2]? r2_3222 : r2_3221;
wire r3_1612;
assign r3_1612 = in[2]? r2_3224 : r2_3223;
wire r3_1613;
assign r3_1613 = in[2]? r2_3226 : r2_3225;
wire r3_1614;
assign r3_1614 = in[2]? r2_3228 : r2_3227;
wire r3_1615;
assign r3_1615 = in[2]? r2_3230 : r2_3229;
wire r3_1616;
assign r3_1616 = in[2]? r2_3232 : r2_3231;
wire r3_1617;
assign r3_1617 = in[2]? r2_3234 : r2_3233;
wire r3_1618;
assign r3_1618 = in[2]? r2_3236 : r2_3235;
wire r3_1619;
assign r3_1619 = in[2]? r2_3238 : r2_3237;
wire r3_1620;
assign r3_1620 = in[2]? r2_3240 : r2_3239;
wire r3_1621;
assign r3_1621 = in[2]? r2_3242 : r2_3241;
wire r3_1622;
assign r3_1622 = in[2]? r2_3244 : r2_3243;
wire r3_1623;
assign r3_1623 = in[2]? r2_3246 : r2_3245;
wire r3_1624;
assign r3_1624 = in[2]? r2_3248 : r2_3247;
wire r3_1625;
assign r3_1625 = in[2]? r2_3250 : r2_3249;
wire r3_1626;
assign r3_1626 = in[2]? r2_3252 : r2_3251;
wire r3_1627;
assign r3_1627 = in[2]? r2_3254 : r2_3253;
wire r3_1628;
assign r3_1628 = in[2]? r2_3256 : r2_3255;
wire r3_1629;
assign r3_1629 = in[2]? r2_3258 : r2_3257;
wire r3_1630;
assign r3_1630 = in[2]? r2_3260 : r2_3259;
wire r3_1631;
assign r3_1631 = in[2]? r2_3262 : r2_3261;
wire r3_1632;
assign r3_1632 = in[2]? r2_3264 : r2_3263;
wire r3_1633;
assign r3_1633 = in[2]? r2_3266 : r2_3265;
wire r3_1634;
assign r3_1634 = in[2]? r2_3268 : r2_3267;
wire r3_1635;
assign r3_1635 = in[2]? r2_3270 : r2_3269;
wire r3_1636;
assign r3_1636 = in[2]? r2_3272 : r2_3271;
wire r3_1637;
assign r3_1637 = in[2]? r2_3274 : r2_3273;
wire r3_1638;
assign r3_1638 = in[2]? r2_3276 : r2_3275;
wire r3_1639;
assign r3_1639 = in[2]? r2_3278 : r2_3277;
wire r3_1640;
assign r3_1640 = in[2]? r2_3280 : r2_3279;
wire r3_1641;
assign r3_1641 = in[2]? r2_3282 : r2_3281;
wire r3_1642;
assign r3_1642 = in[2]? r2_3284 : r2_3283;
wire r3_1643;
assign r3_1643 = in[2]? r2_3286 : r2_3285;
wire r3_1644;
assign r3_1644 = in[2]? r2_3288 : r2_3287;
wire r3_1645;
assign r3_1645 = in[2]? r2_3290 : r2_3289;
wire r3_1646;
assign r3_1646 = in[2]? r2_3292 : r2_3291;
wire r3_1647;
assign r3_1647 = in[2]? r2_3294 : r2_3293;
wire r3_1648;
assign r3_1648 = in[2]? r2_3296 : r2_3295;
wire r3_1649;
assign r3_1649 = in[2]? r2_3298 : r2_3297;
wire r3_1650;
assign r3_1650 = in[2]? r2_3300 : r2_3299;
wire r3_1651;
assign r3_1651 = in[2]? r2_3302 : r2_3301;
wire r3_1652;
assign r3_1652 = in[2]? r2_3304 : r2_3303;
wire r3_1653;
assign r3_1653 = in[2]? r2_3306 : r2_3305;
wire r3_1654;
assign r3_1654 = in[2]? r2_3308 : r2_3307;
wire r3_1655;
assign r3_1655 = in[2]? r2_3310 : r2_3309;
wire r3_1656;
assign r3_1656 = in[2]? r2_3312 : r2_3311;
wire r3_1657;
assign r3_1657 = in[2]? r2_3314 : r2_3313;
wire r3_1658;
assign r3_1658 = in[2]? r2_3316 : r2_3315;
wire r3_1659;
assign r3_1659 = in[2]? r2_3318 : r2_3317;
wire r3_1660;
assign r3_1660 = in[2]? r2_3320 : r2_3319;
wire r3_1661;
assign r3_1661 = in[2]? r2_3322 : r2_3321;
wire r3_1662;
assign r3_1662 = in[2]? r2_3324 : r2_3323;
wire r3_1663;
assign r3_1663 = in[2]? r2_3326 : r2_3325;
wire r3_1664;
assign r3_1664 = in[2]? r2_3328 : r2_3327;
wire r3_1665;
assign r3_1665 = in[2]? r2_3330 : r2_3329;
wire r3_1666;
assign r3_1666 = in[2]? r2_3332 : r2_3331;
wire r3_1667;
assign r3_1667 = in[2]? r2_3334 : r2_3333;
wire r3_1668;
assign r3_1668 = in[2]? r2_3336 : r2_3335;
wire r3_1669;
assign r3_1669 = in[2]? r2_3338 : r2_3337;
wire r3_1670;
assign r3_1670 = in[2]? r2_3340 : r2_3339;
wire r3_1671;
assign r3_1671 = in[2]? r2_3342 : r2_3341;
wire r3_1672;
assign r3_1672 = in[2]? r2_3344 : r2_3343;
wire r3_1673;
assign r3_1673 = in[2]? r2_3346 : r2_3345;
wire r3_1674;
assign r3_1674 = in[2]? r2_3348 : r2_3347;
wire r3_1675;
assign r3_1675 = in[2]? r2_3350 : r2_3349;
wire r3_1676;
assign r3_1676 = in[2]? r2_3352 : r2_3351;
wire r3_1677;
assign r3_1677 = in[2]? r2_3354 : r2_3353;
wire r3_1678;
assign r3_1678 = in[2]? r2_3356 : r2_3355;
wire r3_1679;
assign r3_1679 = in[2]? r2_3358 : r2_3357;
wire r3_1680;
assign r3_1680 = in[2]? r2_3360 : r2_3359;
wire r3_1681;
assign r3_1681 = in[2]? r2_3362 : r2_3361;
wire r3_1682;
assign r3_1682 = in[2]? r2_3364 : r2_3363;
wire r3_1683;
assign r3_1683 = in[2]? r2_3366 : r2_3365;
wire r3_1684;
assign r3_1684 = in[2]? r2_3368 : r2_3367;
wire r3_1685;
assign r3_1685 = in[2]? r2_3370 : r2_3369;
wire r3_1686;
assign r3_1686 = in[2]? r2_3372 : r2_3371;
wire r3_1687;
assign r3_1687 = in[2]? r2_3374 : r2_3373;
wire r3_1688;
assign r3_1688 = in[2]? r2_3376 : r2_3375;
wire r3_1689;
assign r3_1689 = in[2]? r2_3378 : r2_3377;
wire r3_1690;
assign r3_1690 = in[2]? r2_3380 : r2_3379;
wire r3_1691;
assign r3_1691 = in[2]? r2_3382 : r2_3381;
wire r3_1692;
assign r3_1692 = in[2]? r2_3384 : r2_3383;
wire r3_1693;
assign r3_1693 = in[2]? r2_3386 : r2_3385;
wire r3_1694;
assign r3_1694 = in[2]? r2_3388 : r2_3387;
wire r3_1695;
assign r3_1695 = in[2]? r2_3390 : r2_3389;
wire r3_1696;
assign r3_1696 = in[2]? r2_3392 : r2_3391;
wire r3_1697;
assign r3_1697 = in[2]? r2_3394 : r2_3393;
wire r3_1698;
assign r3_1698 = in[2]? r2_3396 : r2_3395;
wire r3_1699;
assign r3_1699 = in[2]? r2_3398 : r2_3397;
wire r3_1700;
assign r3_1700 = in[2]? r2_3400 : r2_3399;
wire r3_1701;
assign r3_1701 = in[2]? r2_3402 : r2_3401;
wire r3_1702;
assign r3_1702 = in[2]? r2_3404 : r2_3403;
wire r3_1703;
assign r3_1703 = in[2]? r2_3406 : r2_3405;
wire r3_1704;
assign r3_1704 = in[2]? r2_3408 : r2_3407;
wire r3_1705;
assign r3_1705 = in[2]? r2_3410 : r2_3409;
wire r3_1706;
assign r3_1706 = in[2]? r2_3412 : r2_3411;
wire r3_1707;
assign r3_1707 = in[2]? r2_3414 : r2_3413;
wire r3_1708;
assign r3_1708 = in[2]? r2_3416 : r2_3415;
wire r3_1709;
assign r3_1709 = in[2]? r2_3418 : r2_3417;
wire r3_1710;
assign r3_1710 = in[2]? r2_3420 : r2_3419;
wire r3_1711;
assign r3_1711 = in[2]? r2_3422 : r2_3421;
wire r3_1712;
assign r3_1712 = in[2]? r2_3424 : r2_3423;
wire r3_1713;
assign r3_1713 = in[2]? r2_3426 : r2_3425;
wire r3_1714;
assign r3_1714 = in[2]? r2_3428 : r2_3427;
wire r3_1715;
assign r3_1715 = in[2]? r2_3430 : r2_3429;
wire r3_1716;
assign r3_1716 = in[2]? r2_3432 : r2_3431;
wire r3_1717;
assign r3_1717 = in[2]? r2_3434 : r2_3433;
wire r3_1718;
assign r3_1718 = in[2]? r2_3436 : r2_3435;
wire r3_1719;
assign r3_1719 = in[2]? r2_3438 : r2_3437;
wire r3_1720;
assign r3_1720 = in[2]? r2_3440 : r2_3439;
wire r3_1721;
assign r3_1721 = in[2]? r2_3442 : r2_3441;
wire r3_1722;
assign r3_1722 = in[2]? r2_3444 : r2_3443;
wire r3_1723;
assign r3_1723 = in[2]? r2_3446 : r2_3445;
wire r3_1724;
assign r3_1724 = in[2]? r2_3448 : r2_3447;
wire r3_1725;
assign r3_1725 = in[2]? r2_3450 : r2_3449;
wire r3_1726;
assign r3_1726 = in[2]? r2_3452 : r2_3451;
wire r3_1727;
assign r3_1727 = in[2]? r2_3454 : r2_3453;
wire r3_1728;
assign r3_1728 = in[2]? r2_3456 : r2_3455;
wire r3_1729;
assign r3_1729 = in[2]? r2_3458 : r2_3457;
wire r3_1730;
assign r3_1730 = in[2]? r2_3460 : r2_3459;
wire r3_1731;
assign r3_1731 = in[2]? r2_3462 : r2_3461;
wire r3_1732;
assign r3_1732 = in[2]? r2_3464 : r2_3463;
wire r3_1733;
assign r3_1733 = in[2]? r2_3466 : r2_3465;
wire r3_1734;
assign r3_1734 = in[2]? r2_3468 : r2_3467;
wire r3_1735;
assign r3_1735 = in[2]? r2_3470 : r2_3469;
wire r3_1736;
assign r3_1736 = in[2]? r2_3472 : r2_3471;
wire r3_1737;
assign r3_1737 = in[2]? r2_3474 : r2_3473;
wire r3_1738;
assign r3_1738 = in[2]? r2_3476 : r2_3475;
wire r3_1739;
assign r3_1739 = in[2]? r2_3478 : r2_3477;
wire r3_1740;
assign r3_1740 = in[2]? r2_3480 : r2_3479;
wire r3_1741;
assign r3_1741 = in[2]? r2_3482 : r2_3481;
wire r3_1742;
assign r3_1742 = in[2]? r2_3484 : r2_3483;
wire r3_1743;
assign r3_1743 = in[2]? r2_3486 : r2_3485;
wire r3_1744;
assign r3_1744 = in[2]? r2_3488 : r2_3487;
wire r3_1745;
assign r3_1745 = in[2]? r2_3490 : r2_3489;
wire r3_1746;
assign r3_1746 = in[2]? r2_3492 : r2_3491;
wire r3_1747;
assign r3_1747 = in[2]? r2_3494 : r2_3493;
wire r3_1748;
assign r3_1748 = in[2]? r2_3496 : r2_3495;
wire r3_1749;
assign r3_1749 = in[2]? r2_3498 : r2_3497;
wire r3_1750;
assign r3_1750 = in[2]? r2_3500 : r2_3499;
wire r3_1751;
assign r3_1751 = in[2]? r2_3502 : r2_3501;
wire r3_1752;
assign r3_1752 = in[2]? r2_3504 : r2_3503;
wire r3_1753;
assign r3_1753 = in[2]? r2_3506 : r2_3505;
wire r3_1754;
assign r3_1754 = in[2]? r2_3508 : r2_3507;
wire r3_1755;
assign r3_1755 = in[2]? r2_3510 : r2_3509;
wire r3_1756;
assign r3_1756 = in[2]? r2_3512 : r2_3511;
wire r3_1757;
assign r3_1757 = in[2]? r2_3514 : r2_3513;
wire r3_1758;
assign r3_1758 = in[2]? r2_3516 : r2_3515;
wire r3_1759;
assign r3_1759 = in[2]? r2_3518 : r2_3517;
wire r3_1760;
assign r3_1760 = in[2]? r2_3520 : r2_3519;
wire r3_1761;
assign r3_1761 = in[2]? r2_3522 : r2_3521;
wire r3_1762;
assign r3_1762 = in[2]? r2_3524 : r2_3523;
wire r3_1763;
assign r3_1763 = in[2]? r2_3526 : r2_3525;
wire r3_1764;
assign r3_1764 = in[2]? r2_3528 : r2_3527;
wire r3_1765;
assign r3_1765 = in[2]? r2_3530 : r2_3529;
wire r3_1766;
assign r3_1766 = in[2]? r2_3532 : r2_3531;
wire r3_1767;
assign r3_1767 = in[2]? r2_3534 : r2_3533;
wire r3_1768;
assign r3_1768 = in[2]? r2_3536 : r2_3535;
wire r3_1769;
assign r3_1769 = in[2]? r2_3538 : r2_3537;
wire r3_1770;
assign r3_1770 = in[2]? r2_3540 : r2_3539;
wire r3_1771;
assign r3_1771 = in[2]? r2_3542 : r2_3541;
wire r3_1772;
assign r3_1772 = in[2]? r2_3544 : r2_3543;
wire r3_1773;
assign r3_1773 = in[2]? r2_3546 : r2_3545;
wire r3_1774;
assign r3_1774 = in[2]? r2_3548 : r2_3547;
wire r3_1775;
assign r3_1775 = in[2]? r2_3550 : r2_3549;
wire r3_1776;
assign r3_1776 = in[2]? r2_3552 : r2_3551;
wire r3_1777;
assign r3_1777 = in[2]? r2_3554 : r2_3553;
wire r3_1778;
assign r3_1778 = in[2]? r2_3556 : r2_3555;
wire r3_1779;
assign r3_1779 = in[2]? r2_3558 : r2_3557;
wire r3_1780;
assign r3_1780 = in[2]? r2_3560 : r2_3559;
wire r3_1781;
assign r3_1781 = in[2]? r2_3562 : r2_3561;
wire r3_1782;
assign r3_1782 = in[2]? r2_3564 : r2_3563;
wire r3_1783;
assign r3_1783 = in[2]? r2_3566 : r2_3565;
wire r3_1784;
assign r3_1784 = in[2]? r2_3568 : r2_3567;
wire r3_1785;
assign r3_1785 = in[2]? r2_3570 : r2_3569;
wire r3_1786;
assign r3_1786 = in[2]? r2_3572 : r2_3571;
wire r3_1787;
assign r3_1787 = in[2]? r2_3574 : r2_3573;
wire r3_1788;
assign r3_1788 = in[2]? r2_3576 : r2_3575;
wire r3_1789;
assign r3_1789 = in[2]? r2_3578 : r2_3577;
wire r3_1790;
assign r3_1790 = in[2]? r2_3580 : r2_3579;
wire r3_1791;
assign r3_1791 = in[2]? r2_3582 : r2_3581;
wire r3_1792;
assign r3_1792 = in[2]? r2_3584 : r2_3583;
wire r3_1793;
assign r3_1793 = in[2]? r2_3586 : r2_3585;
wire r3_1794;
assign r3_1794 = in[2]? r2_3588 : r2_3587;
wire r3_1795;
assign r3_1795 = in[2]? r2_3590 : r2_3589;
wire r3_1796;
assign r3_1796 = in[2]? r2_3592 : r2_3591;
wire r3_1797;
assign r3_1797 = in[2]? r2_3594 : r2_3593;
wire r3_1798;
assign r3_1798 = in[2]? r2_3596 : r2_3595;
wire r3_1799;
assign r3_1799 = in[2]? r2_3598 : r2_3597;
wire r3_1800;
assign r3_1800 = in[2]? r2_3600 : r2_3599;
wire r3_1801;
assign r3_1801 = in[2]? r2_3602 : r2_3601;
wire r3_1802;
assign r3_1802 = in[2]? r2_3604 : r2_3603;
wire r3_1803;
assign r3_1803 = in[2]? r2_3606 : r2_3605;
wire r3_1804;
assign r3_1804 = in[2]? r2_3608 : r2_3607;
wire r3_1805;
assign r3_1805 = in[2]? r2_3610 : r2_3609;
wire r3_1806;
assign r3_1806 = in[2]? r2_3612 : r2_3611;
wire r3_1807;
assign r3_1807 = in[2]? r2_3614 : r2_3613;
wire r3_1808;
assign r3_1808 = in[2]? r2_3616 : r2_3615;
wire r3_1809;
assign r3_1809 = in[2]? r2_3618 : r2_3617;
wire r3_1810;
assign r3_1810 = in[2]? r2_3620 : r2_3619;
wire r3_1811;
assign r3_1811 = in[2]? r2_3622 : r2_3621;
wire r3_1812;
assign r3_1812 = in[2]? r2_3624 : r2_3623;
wire r3_1813;
assign r3_1813 = in[2]? r2_3626 : r2_3625;
wire r3_1814;
assign r3_1814 = in[2]? r2_3628 : r2_3627;
wire r3_1815;
assign r3_1815 = in[2]? r2_3630 : r2_3629;
wire r3_1816;
assign r3_1816 = in[2]? r2_3632 : r2_3631;
wire r3_1817;
assign r3_1817 = in[2]? r2_3634 : r2_3633;
wire r3_1818;
assign r3_1818 = in[2]? r2_3636 : r2_3635;
wire r3_1819;
assign r3_1819 = in[2]? r2_3638 : r2_3637;
wire r3_1820;
assign r3_1820 = in[2]? r2_3640 : r2_3639;
wire r3_1821;
assign r3_1821 = in[2]? r2_3642 : r2_3641;
wire r3_1822;
assign r3_1822 = in[2]? r2_3644 : r2_3643;
wire r3_1823;
assign r3_1823 = in[2]? r2_3646 : r2_3645;
wire r3_1824;
assign r3_1824 = in[2]? r2_3648 : r2_3647;
wire r3_1825;
assign r3_1825 = in[2]? r2_3650 : r2_3649;
wire r3_1826;
assign r3_1826 = in[2]? r2_3652 : r2_3651;
wire r3_1827;
assign r3_1827 = in[2]? r2_3654 : r2_3653;
wire r3_1828;
assign r3_1828 = in[2]? r2_3656 : r2_3655;
wire r3_1829;
assign r3_1829 = in[2]? r2_3658 : r2_3657;
wire r3_1830;
assign r3_1830 = in[2]? r2_3660 : r2_3659;
wire r3_1831;
assign r3_1831 = in[2]? r2_3662 : r2_3661;
wire r3_1832;
assign r3_1832 = in[2]? r2_3664 : r2_3663;
wire r3_1833;
assign r3_1833 = in[2]? r2_3666 : r2_3665;
wire r3_1834;
assign r3_1834 = in[2]? r2_3668 : r2_3667;
wire r3_1835;
assign r3_1835 = in[2]? r2_3670 : r2_3669;
wire r3_1836;
assign r3_1836 = in[2]? r2_3672 : r2_3671;
wire r3_1837;
assign r3_1837 = in[2]? r2_3674 : r2_3673;
wire r3_1838;
assign r3_1838 = in[2]? r2_3676 : r2_3675;
wire r3_1839;
assign r3_1839 = in[2]? r2_3678 : r2_3677;
wire r3_1840;
assign r3_1840 = in[2]? r2_3680 : r2_3679;
wire r3_1841;
assign r3_1841 = in[2]? r2_3682 : r2_3681;
wire r3_1842;
assign r3_1842 = in[2]? r2_3684 : r2_3683;
wire r3_1843;
assign r3_1843 = in[2]? r2_3686 : r2_3685;
wire r3_1844;
assign r3_1844 = in[2]? r2_3688 : r2_3687;
wire r3_1845;
assign r3_1845 = in[2]? r2_3690 : r2_3689;
wire r3_1846;
assign r3_1846 = in[2]? r2_3692 : r2_3691;
wire r3_1847;
assign r3_1847 = in[2]? r2_3694 : r2_3693;
wire r3_1848;
assign r3_1848 = in[2]? r2_3696 : r2_3695;
wire r3_1849;
assign r3_1849 = in[2]? r2_3698 : r2_3697;
wire r3_1850;
assign r3_1850 = in[2]? r2_3700 : r2_3699;
wire r3_1851;
assign r3_1851 = in[2]? r2_3702 : r2_3701;
wire r3_1852;
assign r3_1852 = in[2]? r2_3704 : r2_3703;
wire r3_1853;
assign r3_1853 = in[2]? r2_3706 : r2_3705;
wire r3_1854;
assign r3_1854 = in[2]? r2_3708 : r2_3707;
wire r3_1855;
assign r3_1855 = in[2]? r2_3710 : r2_3709;
wire r3_1856;
assign r3_1856 = in[2]? r2_3712 : r2_3711;
wire r3_1857;
assign r3_1857 = in[2]? r2_3714 : r2_3713;
wire r3_1858;
assign r3_1858 = in[2]? r2_3716 : r2_3715;
wire r3_1859;
assign r3_1859 = in[2]? r2_3718 : r2_3717;
wire r3_1860;
assign r3_1860 = in[2]? r2_3720 : r2_3719;
wire r3_1861;
assign r3_1861 = in[2]? r2_3722 : r2_3721;
wire r3_1862;
assign r3_1862 = in[2]? r2_3724 : r2_3723;
wire r3_1863;
assign r3_1863 = in[2]? r2_3726 : r2_3725;
wire r3_1864;
assign r3_1864 = in[2]? r2_3728 : r2_3727;
wire r3_1865;
assign r3_1865 = in[2]? r2_3730 : r2_3729;
wire r3_1866;
assign r3_1866 = in[2]? r2_3732 : r2_3731;
wire r3_1867;
assign r3_1867 = in[2]? r2_3734 : r2_3733;
wire r3_1868;
assign r3_1868 = in[2]? r2_3736 : r2_3735;
wire r3_1869;
assign r3_1869 = in[2]? r2_3738 : r2_3737;
wire r3_1870;
assign r3_1870 = in[2]? r2_3740 : r2_3739;
wire r3_1871;
assign r3_1871 = in[2]? r2_3742 : r2_3741;
wire r3_1872;
assign r3_1872 = in[2]? r2_3744 : r2_3743;
wire r3_1873;
assign r3_1873 = in[2]? r2_3746 : r2_3745;
wire r3_1874;
assign r3_1874 = in[2]? r2_3748 : r2_3747;
wire r3_1875;
assign r3_1875 = in[2]? r2_3750 : r2_3749;
wire r3_1876;
assign r3_1876 = in[2]? r2_3752 : r2_3751;
wire r3_1877;
assign r3_1877 = in[2]? r2_3754 : r2_3753;
wire r3_1878;
assign r3_1878 = in[2]? r2_3756 : r2_3755;
wire r3_1879;
assign r3_1879 = in[2]? r2_3758 : r2_3757;
wire r3_1880;
assign r3_1880 = in[2]? r2_3760 : r2_3759;
wire r3_1881;
assign r3_1881 = in[2]? r2_3762 : r2_3761;
wire r3_1882;
assign r3_1882 = in[2]? r2_3764 : r2_3763;
wire r3_1883;
assign r3_1883 = in[2]? r2_3766 : r2_3765;
wire r3_1884;
assign r3_1884 = in[2]? r2_3768 : r2_3767;
wire r3_1885;
assign r3_1885 = in[2]? r2_3770 : r2_3769;
wire r3_1886;
assign r3_1886 = in[2]? r2_3772 : r2_3771;
wire r3_1887;
assign r3_1887 = in[2]? r2_3774 : r2_3773;
wire r3_1888;
assign r3_1888 = in[2]? r2_3776 : r2_3775;
wire r3_1889;
assign r3_1889 = in[2]? r2_3778 : r2_3777;
wire r3_1890;
assign r3_1890 = in[2]? r2_3780 : r2_3779;
wire r3_1891;
assign r3_1891 = in[2]? r2_3782 : r2_3781;
wire r3_1892;
assign r3_1892 = in[2]? r2_3784 : r2_3783;
wire r3_1893;
assign r3_1893 = in[2]? r2_3786 : r2_3785;
wire r3_1894;
assign r3_1894 = in[2]? r2_3788 : r2_3787;
wire r3_1895;
assign r3_1895 = in[2]? r2_3790 : r2_3789;
wire r3_1896;
assign r3_1896 = in[2]? r2_3792 : r2_3791;
wire r3_1897;
assign r3_1897 = in[2]? r2_3794 : r2_3793;
wire r3_1898;
assign r3_1898 = in[2]? r2_3796 : r2_3795;
wire r3_1899;
assign r3_1899 = in[2]? r2_3798 : r2_3797;
wire r3_1900;
assign r3_1900 = in[2]? r2_3800 : r2_3799;
wire r3_1901;
assign r3_1901 = in[2]? r2_3802 : r2_3801;
wire r3_1902;
assign r3_1902 = in[2]? r2_3804 : r2_3803;
wire r3_1903;
assign r3_1903 = in[2]? r2_3806 : r2_3805;
wire r3_1904;
assign r3_1904 = in[2]? r2_3808 : r2_3807;
wire r3_1905;
assign r3_1905 = in[2]? r2_3810 : r2_3809;
wire r3_1906;
assign r3_1906 = in[2]? r2_3812 : r2_3811;
wire r3_1907;
assign r3_1907 = in[2]? r2_3814 : r2_3813;
wire r3_1908;
assign r3_1908 = in[2]? r2_3816 : r2_3815;
wire r3_1909;
assign r3_1909 = in[2]? r2_3818 : r2_3817;
wire r3_1910;
assign r3_1910 = in[2]? r2_3820 : r2_3819;
wire r3_1911;
assign r3_1911 = in[2]? r2_3822 : r2_3821;
wire r3_1912;
assign r3_1912 = in[2]? r2_3824 : r2_3823;
wire r3_1913;
assign r3_1913 = in[2]? r2_3826 : r2_3825;
wire r3_1914;
assign r3_1914 = in[2]? r2_3828 : r2_3827;
wire r3_1915;
assign r3_1915 = in[2]? r2_3830 : r2_3829;
wire r3_1916;
assign r3_1916 = in[2]? r2_3832 : r2_3831;
wire r3_1917;
assign r3_1917 = in[2]? r2_3834 : r2_3833;
wire r3_1918;
assign r3_1918 = in[2]? r2_3836 : r2_3835;
wire r3_1919;
assign r3_1919 = in[2]? r2_3838 : r2_3837;
wire r3_1920;
assign r3_1920 = in[2]? r2_3840 : r2_3839;
wire r3_1921;
assign r3_1921 = in[2]? r2_3842 : r2_3841;
wire r3_1922;
assign r3_1922 = in[2]? r2_3844 : r2_3843;
wire r3_1923;
assign r3_1923 = in[2]? r2_3846 : r2_3845;
wire r3_1924;
assign r3_1924 = in[2]? r2_3848 : r2_3847;
wire r3_1925;
assign r3_1925 = in[2]? r2_3850 : r2_3849;
wire r3_1926;
assign r3_1926 = in[2]? r2_3852 : r2_3851;
wire r3_1927;
assign r3_1927 = in[2]? r2_3854 : r2_3853;
wire r3_1928;
assign r3_1928 = in[2]? r2_3856 : r2_3855;
wire r3_1929;
assign r3_1929 = in[2]? r2_3858 : r2_3857;
wire r3_1930;
assign r3_1930 = in[2]? r2_3860 : r2_3859;
wire r3_1931;
assign r3_1931 = in[2]? r2_3862 : r2_3861;
wire r3_1932;
assign r3_1932 = in[2]? r2_3864 : r2_3863;
wire r3_1933;
assign r3_1933 = in[2]? r2_3866 : r2_3865;
wire r3_1934;
assign r3_1934 = in[2]? r2_3868 : r2_3867;
wire r3_1935;
assign r3_1935 = in[2]? r2_3870 : r2_3869;
wire r3_1936;
assign r3_1936 = in[2]? r2_3872 : r2_3871;
wire r3_1937;
assign r3_1937 = in[2]? r2_3874 : r2_3873;
wire r3_1938;
assign r3_1938 = in[2]? r2_3876 : r2_3875;
wire r3_1939;
assign r3_1939 = in[2]? r2_3878 : r2_3877;
wire r3_1940;
assign r3_1940 = in[2]? r2_3880 : r2_3879;
wire r3_1941;
assign r3_1941 = in[2]? r2_3882 : r2_3881;
wire r3_1942;
assign r3_1942 = in[2]? r2_3884 : r2_3883;
wire r3_1943;
assign r3_1943 = in[2]? r2_3886 : r2_3885;
wire r3_1944;
assign r3_1944 = in[2]? r2_3888 : r2_3887;
wire r3_1945;
assign r3_1945 = in[2]? r2_3890 : r2_3889;
wire r3_1946;
assign r3_1946 = in[2]? r2_3892 : r2_3891;
wire r3_1947;
assign r3_1947 = in[2]? r2_3894 : r2_3893;
wire r3_1948;
assign r3_1948 = in[2]? r2_3896 : r2_3895;
wire r3_1949;
assign r3_1949 = in[2]? r2_3898 : r2_3897;
wire r3_1950;
assign r3_1950 = in[2]? r2_3900 : r2_3899;
wire r3_1951;
assign r3_1951 = in[2]? r2_3902 : r2_3901;
wire r3_1952;
assign r3_1952 = in[2]? r2_3904 : r2_3903;
wire r3_1953;
assign r3_1953 = in[2]? r2_3906 : r2_3905;
wire r3_1954;
assign r3_1954 = in[2]? r2_3908 : r2_3907;
wire r3_1955;
assign r3_1955 = in[2]? r2_3910 : r2_3909;
wire r3_1956;
assign r3_1956 = in[2]? r2_3912 : r2_3911;
wire r3_1957;
assign r3_1957 = in[2]? r2_3914 : r2_3913;
wire r3_1958;
assign r3_1958 = in[2]? r2_3916 : r2_3915;
wire r3_1959;
assign r3_1959 = in[2]? r2_3918 : r2_3917;
wire r3_1960;
assign r3_1960 = in[2]? r2_3920 : r2_3919;
wire r3_1961;
assign r3_1961 = in[2]? r2_3922 : r2_3921;
wire r3_1962;
assign r3_1962 = in[2]? r2_3924 : r2_3923;
wire r3_1963;
assign r3_1963 = in[2]? r2_3926 : r2_3925;
wire r3_1964;
assign r3_1964 = in[2]? r2_3928 : r2_3927;
wire r3_1965;
assign r3_1965 = in[2]? r2_3930 : r2_3929;
wire r3_1966;
assign r3_1966 = in[2]? r2_3932 : r2_3931;
wire r3_1967;
assign r3_1967 = in[2]? r2_3934 : r2_3933;
wire r3_1968;
assign r3_1968 = in[2]? r2_3936 : r2_3935;
wire r3_1969;
assign r3_1969 = in[2]? r2_3938 : r2_3937;
wire r3_1970;
assign r3_1970 = in[2]? r2_3940 : r2_3939;
wire r3_1971;
assign r3_1971 = in[2]? r2_3942 : r2_3941;
wire r3_1972;
assign r3_1972 = in[2]? r2_3944 : r2_3943;
wire r3_1973;
assign r3_1973 = in[2]? r2_3946 : r2_3945;
wire r3_1974;
assign r3_1974 = in[2]? r2_3948 : r2_3947;
wire r3_1975;
assign r3_1975 = in[2]? r2_3950 : r2_3949;
wire r3_1976;
assign r3_1976 = in[2]? r2_3952 : r2_3951;
wire r3_1977;
assign r3_1977 = in[2]? r2_3954 : r2_3953;
wire r3_1978;
assign r3_1978 = in[2]? r2_3956 : r2_3955;
wire r3_1979;
assign r3_1979 = in[2]? r2_3958 : r2_3957;
wire r3_1980;
assign r3_1980 = in[2]? r2_3960 : r2_3959;
wire r3_1981;
assign r3_1981 = in[2]? r2_3962 : r2_3961;
wire r3_1982;
assign r3_1982 = in[2]? r2_3964 : r2_3963;
wire r3_1983;
assign r3_1983 = in[2]? r2_3966 : r2_3965;
wire r3_1984;
assign r3_1984 = in[2]? r2_3968 : r2_3967;
wire r3_1985;
assign r3_1985 = in[2]? r2_3970 : r2_3969;
wire r3_1986;
assign r3_1986 = in[2]? r2_3972 : r2_3971;
wire r3_1987;
assign r3_1987 = in[2]? r2_3974 : r2_3973;
wire r3_1988;
assign r3_1988 = in[2]? r2_3976 : r2_3975;
wire r3_1989;
assign r3_1989 = in[2]? r2_3978 : r2_3977;
wire r3_1990;
assign r3_1990 = in[2]? r2_3980 : r2_3979;
wire r3_1991;
assign r3_1991 = in[2]? r2_3982 : r2_3981;
wire r3_1992;
assign r3_1992 = in[2]? r2_3984 : r2_3983;
wire r3_1993;
assign r3_1993 = in[2]? r2_3986 : r2_3985;
wire r3_1994;
assign r3_1994 = in[2]? r2_3988 : r2_3987;
wire r3_1995;
assign r3_1995 = in[2]? r2_3990 : r2_3989;
wire r3_1996;
assign r3_1996 = in[2]? r2_3992 : r2_3991;
wire r3_1997;
assign r3_1997 = in[2]? r2_3994 : r2_3993;
wire r3_1998;
assign r3_1998 = in[2]? r2_3996 : r2_3995;
wire r3_1999;
assign r3_1999 = in[2]? r2_3998 : r2_3997;
wire r3_2000;
assign r3_2000 = in[2]? r2_4000 : r2_3999;
wire r3_2001;
assign r3_2001 = in[2]? r2_4002 : r2_4001;
wire r3_2002;
assign r3_2002 = in[2]? r2_4004 : r2_4003;
wire r3_2003;
assign r3_2003 = in[2]? r2_4006 : r2_4005;
wire r3_2004;
assign r3_2004 = in[2]? r2_4008 : r2_4007;
wire r3_2005;
assign r3_2005 = in[2]? r2_4010 : r2_4009;
wire r3_2006;
assign r3_2006 = in[2]? r2_4012 : r2_4011;
wire r3_2007;
assign r3_2007 = in[2]? r2_4014 : r2_4013;
wire r3_2008;
assign r3_2008 = in[2]? r2_4016 : r2_4015;
wire r3_2009;
assign r3_2009 = in[2]? r2_4018 : r2_4017;
wire r3_2010;
assign r3_2010 = in[2]? r2_4020 : r2_4019;
wire r3_2011;
assign r3_2011 = in[2]? r2_4022 : r2_4021;
wire r3_2012;
assign r3_2012 = in[2]? r2_4024 : r2_4023;
wire r3_2013;
assign r3_2013 = in[2]? r2_4026 : r2_4025;
wire r3_2014;
assign r3_2014 = in[2]? r2_4028 : r2_4027;
wire r3_2015;
assign r3_2015 = in[2]? r2_4030 : r2_4029;
wire r3_2016;
assign r3_2016 = in[2]? r2_4032 : r2_4031;
wire r3_2017;
assign r3_2017 = in[2]? r2_4034 : r2_4033;
wire r3_2018;
assign r3_2018 = in[2]? r2_4036 : r2_4035;
wire r3_2019;
assign r3_2019 = in[2]? r2_4038 : r2_4037;
wire r3_2020;
assign r3_2020 = in[2]? r2_4040 : r2_4039;
wire r3_2021;
assign r3_2021 = in[2]? r2_4042 : r2_4041;
wire r3_2022;
assign r3_2022 = in[2]? r2_4044 : r2_4043;
wire r3_2023;
assign r3_2023 = in[2]? r2_4046 : r2_4045;
wire r3_2024;
assign r3_2024 = in[2]? r2_4048 : r2_4047;
wire r3_2025;
assign r3_2025 = in[2]? r2_4050 : r2_4049;
wire r3_2026;
assign r3_2026 = in[2]? r2_4052 : r2_4051;
wire r3_2027;
assign r3_2027 = in[2]? r2_4054 : r2_4053;
wire r3_2028;
assign r3_2028 = in[2]? r2_4056 : r2_4055;
wire r3_2029;
assign r3_2029 = in[2]? r2_4058 : r2_4057;
wire r3_2030;
assign r3_2030 = in[2]? r2_4060 : r2_4059;
wire r3_2031;
assign r3_2031 = in[2]? r2_4062 : r2_4061;
wire r3_2032;
assign r3_2032 = in[2]? r2_4064 : r2_4063;
wire r3_2033;
assign r3_2033 = in[2]? r2_4066 : r2_4065;
wire r3_2034;
assign r3_2034 = in[2]? r2_4068 : r2_4067;
wire r3_2035;
assign r3_2035 = in[2]? r2_4070 : r2_4069;
wire r3_2036;
assign r3_2036 = in[2]? r2_4072 : r2_4071;
wire r3_2037;
assign r3_2037 = in[2]? r2_4074 : r2_4073;
wire r3_2038;
assign r3_2038 = in[2]? r2_4076 : r2_4075;
wire r3_2039;
assign r3_2039 = in[2]? r2_4078 : r2_4077;
wire r3_2040;
assign r3_2040 = in[2]? r2_4080 : r2_4079;
wire r3_2041;
assign r3_2041 = in[2]? r2_4082 : r2_4081;
wire r3_2042;
assign r3_2042 = in[2]? r2_4084 : r2_4083;
wire r3_2043;
assign r3_2043 = in[2]? r2_4086 : r2_4085;
wire r3_2044;
assign r3_2044 = in[2]? r2_4088 : r2_4087;
wire r3_2045;
assign r3_2045 = in[2]? r2_4090 : r2_4089;
wire r3_2046;
assign r3_2046 = in[2]? r2_4092 : r2_4091;
wire r3_2047;
assign r3_2047 = in[2]? r2_4094 : r2_4093;
wire r3_2048;
assign r3_2048 = in[2]? r2_4096 : r2_4095;
wire r3_2049;
assign r3_2049 = in[2]? r2_4098 : r2_4097;
wire r3_2050;
assign r3_2050 = in[2]? r2_4100 : r2_4099;
wire r3_2051;
assign r3_2051 = in[2]? r2_4102 : r2_4101;
wire r3_2052;
assign r3_2052 = in[2]? r2_4104 : r2_4103;
wire r3_2053;
assign r3_2053 = in[2]? r2_4106 : r2_4105;
wire r3_2054;
assign r3_2054 = in[2]? r2_4108 : r2_4107;
wire r3_2055;
assign r3_2055 = in[2]? r2_4110 : r2_4109;
wire r3_2056;
assign r3_2056 = in[2]? r2_4112 : r2_4111;
wire r3_2057;
assign r3_2057 = in[2]? r2_4114 : r2_4113;
wire r3_2058;
assign r3_2058 = in[2]? r2_4116 : r2_4115;
wire r3_2059;
assign r3_2059 = in[2]? r2_4118 : r2_4117;
wire r3_2060;
assign r3_2060 = in[2]? r2_4120 : r2_4119;
wire r3_2061;
assign r3_2061 = in[2]? r2_4122 : r2_4121;
wire r3_2062;
assign r3_2062 = in[2]? r2_4124 : r2_4123;
wire r3_2063;
assign r3_2063 = in[2]? r2_4126 : r2_4125;
wire r3_2064;
assign r3_2064 = in[2]? r2_4128 : r2_4127;
wire r3_2065;
assign r3_2065 = in[2]? r2_4130 : r2_4129;
wire r3_2066;
assign r3_2066 = in[2]? r2_4132 : r2_4131;
wire r3_2067;
assign r3_2067 = in[2]? r2_4134 : r2_4133;
wire r3_2068;
assign r3_2068 = in[2]? r2_4136 : r2_4135;
wire r3_2069;
assign r3_2069 = in[2]? r2_4138 : r2_4137;
wire r3_2070;
assign r3_2070 = in[2]? r2_4140 : r2_4139;
wire r3_2071;
assign r3_2071 = in[2]? r2_4142 : r2_4141;
wire r3_2072;
assign r3_2072 = in[2]? r2_4144 : r2_4143;
wire r3_2073;
assign r3_2073 = in[2]? r2_4146 : r2_4145;
wire r3_2074;
assign r3_2074 = in[2]? r2_4148 : r2_4147;
wire r3_2075;
assign r3_2075 = in[2]? r2_4150 : r2_4149;
wire r3_2076;
assign r3_2076 = in[2]? r2_4152 : r2_4151;
wire r3_2077;
assign r3_2077 = in[2]? r2_4154 : r2_4153;
wire r3_2078;
assign r3_2078 = in[2]? r2_4156 : r2_4155;
wire r3_2079;
assign r3_2079 = in[2]? r2_4158 : r2_4157;
wire r3_2080;
assign r3_2080 = in[2]? r2_4160 : r2_4159;
wire r3_2081;
assign r3_2081 = in[2]? r2_4162 : r2_4161;
wire r3_2082;
assign r3_2082 = in[2]? r2_4164 : r2_4163;
wire r3_2083;
assign r3_2083 = in[2]? r2_4166 : r2_4165;
wire r3_2084;
assign r3_2084 = in[2]? r2_4168 : r2_4167;
wire r3_2085;
assign r3_2085 = in[2]? r2_4170 : r2_4169;
wire r3_2086;
assign r3_2086 = in[2]? r2_4172 : r2_4171;
wire r3_2087;
assign r3_2087 = in[2]? r2_4174 : r2_4173;
wire r3_2088;
assign r3_2088 = in[2]? r2_4176 : r2_4175;
wire r3_2089;
assign r3_2089 = in[2]? r2_4178 : r2_4177;
wire r3_2090;
assign r3_2090 = in[2]? r2_4180 : r2_4179;
wire r3_2091;
assign r3_2091 = in[2]? r2_4182 : r2_4181;
wire r3_2092;
assign r3_2092 = in[2]? r2_4184 : r2_4183;
wire r3_2093;
assign r3_2093 = in[2]? r2_4186 : r2_4185;
wire r3_2094;
assign r3_2094 = in[2]? r2_4188 : r2_4187;
wire r3_2095;
assign r3_2095 = in[2]? r2_4190 : r2_4189;
wire r3_2096;
assign r3_2096 = in[2]? r2_4192 : r2_4191;
wire r3_2097;
assign r3_2097 = in[2]? r2_4194 : r2_4193;
wire r3_2098;
assign r3_2098 = in[2]? r2_4196 : r2_4195;
wire r3_2099;
assign r3_2099 = in[2]? r2_4198 : r2_4197;
wire r3_2100;
assign r3_2100 = in[2]? r2_4200 : r2_4199;
wire r3_2101;
assign r3_2101 = in[2]? r2_4202 : r2_4201;
wire r3_2102;
assign r3_2102 = in[2]? r2_4204 : r2_4203;
wire r3_2103;
assign r3_2103 = in[2]? r2_4206 : r2_4205;
wire r3_2104;
assign r3_2104 = in[2]? r2_4208 : r2_4207;
wire r3_2105;
assign r3_2105 = in[2]? r2_4210 : r2_4209;
wire r3_2106;
assign r3_2106 = in[2]? r2_4212 : r2_4211;
wire r3_2107;
assign r3_2107 = in[2]? r2_4214 : r2_4213;
wire r3_2108;
assign r3_2108 = in[2]? r2_4216 : r2_4215;
wire r3_2109;
assign r3_2109 = in[2]? r2_4218 : r2_4217;
wire r3_2110;
assign r3_2110 = in[2]? r2_4220 : r2_4219;
wire r3_2111;
assign r3_2111 = in[2]? r2_4222 : r2_4221;
wire r3_2112;
assign r3_2112 = in[2]? r2_4224 : r2_4223;
wire r3_2113;
assign r3_2113 = in[2]? r2_4226 : r2_4225;
wire r3_2114;
assign r3_2114 = in[2]? r2_4228 : r2_4227;
wire r3_2115;
assign r3_2115 = in[2]? r2_4230 : r2_4229;
wire r3_2116;
assign r3_2116 = in[2]? r2_4232 : r2_4231;
wire r3_2117;
assign r3_2117 = in[2]? r2_4234 : r2_4233;
wire r3_2118;
assign r3_2118 = in[2]? r2_4236 : r2_4235;
wire r3_2119;
assign r3_2119 = in[2]? r2_4238 : r2_4237;
wire r3_2120;
assign r3_2120 = in[2]? r2_4240 : r2_4239;
wire r3_2121;
assign r3_2121 = in[2]? r2_4242 : r2_4241;
wire r3_2122;
assign r3_2122 = in[2]? r2_4244 : r2_4243;
wire r3_2123;
assign r3_2123 = in[2]? r2_4246 : r2_4245;
wire r3_2124;
assign r3_2124 = in[2]? r2_4248 : r2_4247;
wire r3_2125;
assign r3_2125 = in[2]? r2_4250 : r2_4249;
wire r3_2126;
assign r3_2126 = in[2]? r2_4252 : r2_4251;
wire r3_2127;
assign r3_2127 = in[2]? r2_4254 : r2_4253;
wire r3_2128;
assign r3_2128 = in[2]? r2_4256 : r2_4255;
wire r3_2129;
assign r3_2129 = in[2]? r2_4258 : r2_4257;
wire r3_2130;
assign r3_2130 = in[2]? r2_4260 : r2_4259;
wire r3_2131;
assign r3_2131 = in[2]? r2_4262 : r2_4261;
wire r3_2132;
assign r3_2132 = in[2]? r2_4264 : r2_4263;
wire r3_2133;
assign r3_2133 = in[2]? r2_4266 : r2_4265;
wire r3_2134;
assign r3_2134 = in[2]? r2_4268 : r2_4267;
wire r3_2135;
assign r3_2135 = in[2]? r2_4270 : r2_4269;
wire r3_2136;
assign r3_2136 = in[2]? r2_4272 : r2_4271;
wire r3_2137;
assign r3_2137 = in[2]? r2_4274 : r2_4273;
wire r3_2138;
assign r3_2138 = in[2]? r2_4276 : r2_4275;
wire r3_2139;
assign r3_2139 = in[2]? r2_4278 : r2_4277;
wire r3_2140;
assign r3_2140 = in[2]? r2_4280 : r2_4279;
wire r3_2141;
assign r3_2141 = in[2]? r2_4282 : r2_4281;
wire r3_2142;
assign r3_2142 = in[2]? r2_4284 : r2_4283;
wire r3_2143;
assign r3_2143 = in[2]? r2_4286 : r2_4285;
wire r3_2144;
assign r3_2144 = in[2]? r2_4288 : r2_4287;
wire r3_2145;
assign r3_2145 = in[2]? r2_4290 : r2_4289;
wire r3_2146;
assign r3_2146 = in[2]? r2_4292 : r2_4291;
wire r3_2147;
assign r3_2147 = in[2]? r2_4294 : r2_4293;
wire r3_2148;
assign r3_2148 = in[2]? r2_4296 : r2_4295;
wire r3_2149;
assign r3_2149 = in[2]? r2_4298 : r2_4297;
wire r3_2150;
assign r3_2150 = in[2]? r2_4300 : r2_4299;
wire r3_2151;
assign r3_2151 = in[2]? r2_4302 : r2_4301;
wire r3_2152;
assign r3_2152 = in[2]? r2_4304 : r2_4303;
wire r3_2153;
assign r3_2153 = in[2]? r2_4306 : r2_4305;
wire r3_2154;
assign r3_2154 = in[2]? r2_4308 : r2_4307;
wire r3_2155;
assign r3_2155 = in[2]? r2_4310 : r2_4309;
wire r3_2156;
assign r3_2156 = in[2]? r2_4312 : r2_4311;
wire r3_2157;
assign r3_2157 = in[2]? r2_4314 : r2_4313;
wire r3_2158;
assign r3_2158 = in[2]? r2_4316 : r2_4315;
wire r3_2159;
assign r3_2159 = in[2]? r2_4318 : r2_4317;
wire r3_2160;
assign r3_2160 = in[2]? r2_4320 : r2_4319;
wire r3_2161;
assign r3_2161 = in[2]? r2_4322 : r2_4321;
wire r3_2162;
assign r3_2162 = in[2]? r2_4324 : r2_4323;
wire r3_2163;
assign r3_2163 = in[2]? r2_4326 : r2_4325;
wire r3_2164;
assign r3_2164 = in[2]? r2_4328 : r2_4327;
wire r3_2165;
assign r3_2165 = in[2]? r2_4330 : r2_4329;
wire r3_2166;
assign r3_2166 = in[2]? r2_4332 : r2_4331;
wire r3_2167;
assign r3_2167 = in[2]? r2_4334 : r2_4333;
wire r3_2168;
assign r3_2168 = in[2]? r2_4336 : r2_4335;
wire r3_2169;
assign r3_2169 = in[2]? r2_4338 : r2_4337;
wire r3_2170;
assign r3_2170 = in[2]? r2_4340 : r2_4339;
wire r3_2171;
assign r3_2171 = in[2]? r2_4342 : r2_4341;
wire r3_2172;
assign r3_2172 = in[2]? r2_4344 : r2_4343;
wire r3_2173;
assign r3_2173 = in[2]? r2_4346 : r2_4345;
wire r3_2174;
assign r3_2174 = in[2]? r2_4348 : r2_4347;
wire r3_2175;
assign r3_2175 = in[2]? r2_4350 : r2_4349;
wire r3_2176;
assign r3_2176 = in[2]? r2_4352 : r2_4351;
wire r3_2177;
assign r3_2177 = in[2]? r2_4354 : r2_4353;
wire r3_2178;
assign r3_2178 = in[2]? r2_4356 : r2_4355;
wire r3_2179;
assign r3_2179 = in[2]? r2_4358 : r2_4357;
wire r3_2180;
assign r3_2180 = in[2]? r2_4360 : r2_4359;
wire r3_2181;
assign r3_2181 = in[2]? r2_4362 : r2_4361;
wire r3_2182;
assign r3_2182 = in[2]? r2_4364 : r2_4363;
wire r3_2183;
assign r3_2183 = in[2]? r2_4366 : r2_4365;
wire r3_2184;
assign r3_2184 = in[2]? r2_4368 : r2_4367;
wire r3_2185;
assign r3_2185 = in[2]? r2_4370 : r2_4369;
wire r3_2186;
assign r3_2186 = in[2]? r2_4372 : r2_4371;
wire r3_2187;
assign r3_2187 = in[2]? r2_4374 : r2_4373;
wire r3_2188;
assign r3_2188 = in[2]? r2_4376 : r2_4375;
wire r3_2189;
assign r3_2189 = in[2]? r2_4378 : r2_4377;
wire r3_2190;
assign r3_2190 = in[2]? r2_4380 : r2_4379;
wire r3_2191;
assign r3_2191 = in[2]? r2_4382 : r2_4381;
wire r3_2192;
assign r3_2192 = in[2]? r2_4384 : r2_4383;
wire r3_2193;
assign r3_2193 = in[2]? r2_4386 : r2_4385;
wire r3_2194;
assign r3_2194 = in[2]? r2_4388 : r2_4387;
wire r3_2195;
assign r3_2195 = in[2]? r2_4390 : r2_4389;
wire r3_2196;
assign r3_2196 = in[2]? r2_4392 : r2_4391;
wire r3_2197;
assign r3_2197 = in[2]? r2_4394 : r2_4393;
wire r3_2198;
assign r3_2198 = in[2]? r2_4396 : r2_4395;
wire r3_2199;
assign r3_2199 = in[2]? r2_4398 : r2_4397;
wire r3_2200;
assign r3_2200 = in[2]? r2_4400 : r2_4399;
wire r3_2201;
assign r3_2201 = in[2]? r2_4402 : r2_4401;
wire r3_2202;
assign r3_2202 = in[2]? r2_4404 : r2_4403;
wire r3_2203;
assign r3_2203 = in[2]? r2_4406 : r2_4405;
wire r3_2204;
assign r3_2204 = in[2]? r2_4408 : r2_4407;
wire r3_2205;
assign r3_2205 = in[2]? r2_4410 : r2_4409;
wire r3_2206;
assign r3_2206 = in[2]? r2_4412 : r2_4411;
wire r3_2207;
assign r3_2207 = in[2]? r2_4414 : r2_4413;
wire r3_2208;
assign r3_2208 = in[2]? r2_4416 : r2_4415;
wire r3_2209;
assign r3_2209 = in[2]? r2_4418 : r2_4417;
wire r3_2210;
assign r3_2210 = in[2]? r2_4420 : r2_4419;
wire r3_2211;
assign r3_2211 = in[2]? r2_4422 : r2_4421;
wire r3_2212;
assign r3_2212 = in[2]? r2_4424 : r2_4423;
wire r3_2213;
assign r3_2213 = in[2]? r2_4426 : r2_4425;
wire r3_2214;
assign r3_2214 = in[2]? r2_4428 : r2_4427;
wire r3_2215;
assign r3_2215 = in[2]? r2_4430 : r2_4429;
wire r3_2216;
assign r3_2216 = in[2]? r2_4432 : r2_4431;
wire r3_2217;
assign r3_2217 = in[2]? r2_4434 : r2_4433;
wire r3_2218;
assign r3_2218 = in[2]? r2_4436 : r2_4435;
wire r3_2219;
assign r3_2219 = in[2]? r2_4438 : r2_4437;
wire r3_2220;
assign r3_2220 = in[2]? r2_4440 : r2_4439;
wire r3_2221;
assign r3_2221 = in[2]? r2_4442 : r2_4441;
wire r3_2222;
assign r3_2222 = in[2]? r2_4444 : r2_4443;
wire r3_2223;
assign r3_2223 = in[2]? r2_4446 : r2_4445;
wire r3_2224;
assign r3_2224 = in[2]? r2_4448 : r2_4447;
wire r3_2225;
assign r3_2225 = in[2]? r2_4450 : r2_4449;
wire r3_2226;
assign r3_2226 = in[2]? r2_4452 : r2_4451;
wire r3_2227;
assign r3_2227 = in[2]? r2_4454 : r2_4453;
wire r3_2228;
assign r3_2228 = in[2]? r2_4456 : r2_4455;
wire r3_2229;
assign r3_2229 = in[2]? r2_4458 : r2_4457;
wire r3_2230;
assign r3_2230 = in[2]? r2_4460 : r2_4459;
wire r3_2231;
assign r3_2231 = in[2]? r2_4462 : r2_4461;
wire r3_2232;
assign r3_2232 = in[2]? r2_4464 : r2_4463;
wire r3_2233;
assign r3_2233 = in[2]? r2_4466 : r2_4465;
wire r3_2234;
assign r3_2234 = in[2]? r2_4468 : r2_4467;
wire r3_2235;
assign r3_2235 = in[2]? r2_4470 : r2_4469;
wire r3_2236;
assign r3_2236 = in[2]? r2_4472 : r2_4471;
wire r3_2237;
assign r3_2237 = in[2]? r2_4474 : r2_4473;
wire r3_2238;
assign r3_2238 = in[2]? r2_4476 : r2_4475;
wire r3_2239;
assign r3_2239 = in[2]? r2_4478 : r2_4477;
wire r3_2240;
assign r3_2240 = in[2]? r2_4480 : r2_4479;
wire r3_2241;
assign r3_2241 = in[2]? r2_4482 : r2_4481;
wire r3_2242;
assign r3_2242 = in[2]? r2_4484 : r2_4483;
wire r3_2243;
assign r3_2243 = in[2]? r2_4486 : r2_4485;
wire r3_2244;
assign r3_2244 = in[2]? r2_4488 : r2_4487;
wire r3_2245;
assign r3_2245 = in[2]? r2_4490 : r2_4489;
wire r3_2246;
assign r3_2246 = in[2]? r2_4492 : r2_4491;
wire r3_2247;
assign r3_2247 = in[2]? r2_4494 : r2_4493;
wire r3_2248;
assign r3_2248 = in[2]? r2_4496 : r2_4495;
wire r3_2249;
assign r3_2249 = in[2]? r2_4498 : r2_4497;
wire r3_2250;
assign r3_2250 = in[2]? r2_4500 : r2_4499;
wire r3_2251;
assign r3_2251 = in[2]? r2_4502 : r2_4501;
wire r3_2252;
assign r3_2252 = in[2]? r2_4504 : r2_4503;
wire r3_2253;
assign r3_2253 = in[2]? r2_4506 : r2_4505;
wire r3_2254;
assign r3_2254 = in[2]? r2_4508 : r2_4507;
wire r3_2255;
assign r3_2255 = in[2]? r2_4510 : r2_4509;
wire r3_2256;
assign r3_2256 = in[2]? r2_4512 : r2_4511;
wire r3_2257;
assign r3_2257 = in[2]? r2_4514 : r2_4513;
wire r3_2258;
assign r3_2258 = in[2]? r2_4516 : r2_4515;
wire r3_2259;
assign r3_2259 = in[2]? r2_4518 : r2_4517;
wire r3_2260;
assign r3_2260 = in[2]? r2_4520 : r2_4519;
wire r3_2261;
assign r3_2261 = in[2]? r2_4522 : r2_4521;
wire r3_2262;
assign r3_2262 = in[2]? r2_4524 : r2_4523;
wire r3_2263;
assign r3_2263 = in[2]? r2_4526 : r2_4525;
wire r3_2264;
assign r3_2264 = in[2]? r2_4528 : r2_4527;
wire r3_2265;
assign r3_2265 = in[2]? r2_4530 : r2_4529;
wire r3_2266;
assign r3_2266 = in[2]? r2_4532 : r2_4531;
wire r3_2267;
assign r3_2267 = in[2]? r2_4534 : r2_4533;
wire r3_2268;
assign r3_2268 = in[2]? r2_4536 : r2_4535;
wire r3_2269;
assign r3_2269 = in[2]? r2_4538 : r2_4537;
wire r3_2270;
assign r3_2270 = in[2]? r2_4540 : r2_4539;
wire r3_2271;
assign r3_2271 = in[2]? r2_4542 : r2_4541;
wire r3_2272;
assign r3_2272 = in[2]? r2_4544 : r2_4543;
wire r3_2273;
assign r3_2273 = in[2]? r2_4546 : r2_4545;
wire r3_2274;
assign r3_2274 = in[2]? r2_4548 : r2_4547;
wire r3_2275;
assign r3_2275 = in[2]? r2_4550 : r2_4549;
wire r3_2276;
assign r3_2276 = in[2]? r2_4552 : r2_4551;
wire r3_2277;
assign r3_2277 = in[2]? r2_4554 : r2_4553;
wire r3_2278;
assign r3_2278 = in[2]? r2_4556 : r2_4555;
wire r3_2279;
assign r3_2279 = in[2]? r2_4558 : r2_4557;
wire r3_2280;
assign r3_2280 = in[2]? r2_4560 : r2_4559;
wire r3_2281;
assign r3_2281 = in[2]? r2_4562 : r2_4561;
wire r3_2282;
assign r3_2282 = in[2]? r2_4564 : r2_4563;
wire r3_2283;
assign r3_2283 = in[2]? r2_4566 : r2_4565;
wire r3_2284;
assign r3_2284 = in[2]? r2_4568 : r2_4567;
wire r3_2285;
assign r3_2285 = in[2]? r2_4570 : r2_4569;
wire r3_2286;
assign r3_2286 = in[2]? r2_4572 : r2_4571;
wire r3_2287;
assign r3_2287 = in[2]? r2_4574 : r2_4573;
wire r3_2288;
assign r3_2288 = in[2]? r2_4576 : r2_4575;
wire r3_2289;
assign r3_2289 = in[2]? r2_4578 : r2_4577;
wire r3_2290;
assign r3_2290 = in[2]? r2_4580 : r2_4579;
wire r3_2291;
assign r3_2291 = in[2]? r2_4582 : r2_4581;
wire r3_2292;
assign r3_2292 = in[2]? r2_4584 : r2_4583;
wire r3_2293;
assign r3_2293 = in[2]? r2_4586 : r2_4585;
wire r3_2294;
assign r3_2294 = in[2]? r2_4588 : r2_4587;
wire r3_2295;
assign r3_2295 = in[2]? r2_4590 : r2_4589;
wire r3_2296;
assign r3_2296 = in[2]? r2_4592 : r2_4591;
wire r3_2297;
assign r3_2297 = in[2]? r2_4594 : r2_4593;
wire r3_2298;
assign r3_2298 = in[2]? r2_4596 : r2_4595;
wire r3_2299;
assign r3_2299 = in[2]? r2_4598 : r2_4597;
wire r3_2300;
assign r3_2300 = in[2]? r2_4600 : r2_4599;
wire r3_2301;
assign r3_2301 = in[2]? r2_4602 : r2_4601;
wire r3_2302;
assign r3_2302 = in[2]? r2_4604 : r2_4603;
wire r3_2303;
assign r3_2303 = in[2]? r2_4606 : r2_4605;
wire r3_2304;
assign r3_2304 = in[2]? r2_4608 : r2_4607;
wire r3_2305;
assign r3_2305 = in[2]? r2_4610 : r2_4609;
wire r3_2306;
assign r3_2306 = in[2]? r2_4612 : r2_4611;
wire r3_2307;
assign r3_2307 = in[2]? r2_4614 : r2_4613;
wire r3_2308;
assign r3_2308 = in[2]? r2_4616 : r2_4615;
wire r3_2309;
assign r3_2309 = in[2]? r2_4618 : r2_4617;
wire r3_2310;
assign r3_2310 = in[2]? r2_4620 : r2_4619;
wire r3_2311;
assign r3_2311 = in[2]? r2_4622 : r2_4621;
wire r3_2312;
assign r3_2312 = in[2]? r2_4624 : r2_4623;
wire r3_2313;
assign r3_2313 = in[2]? r2_4626 : r2_4625;
wire r3_2314;
assign r3_2314 = in[2]? r2_4628 : r2_4627;
wire r3_2315;
assign r3_2315 = in[2]? r2_4630 : r2_4629;
wire r3_2316;
assign r3_2316 = in[2]? r2_4632 : r2_4631;
wire r3_2317;
assign r3_2317 = in[2]? r2_4634 : r2_4633;
wire r3_2318;
assign r3_2318 = in[2]? r2_4636 : r2_4635;
wire r3_2319;
assign r3_2319 = in[2]? r2_4638 : r2_4637;
wire r3_2320;
assign r3_2320 = in[2]? r2_4640 : r2_4639;
wire r3_2321;
assign r3_2321 = in[2]? r2_4642 : r2_4641;
wire r3_2322;
assign r3_2322 = in[2]? r2_4644 : r2_4643;
wire r3_2323;
assign r3_2323 = in[2]? r2_4646 : r2_4645;
wire r3_2324;
assign r3_2324 = in[2]? r2_4648 : r2_4647;
wire r3_2325;
assign r3_2325 = in[2]? r2_4650 : r2_4649;
wire r3_2326;
assign r3_2326 = in[2]? r2_4652 : r2_4651;
wire r3_2327;
assign r3_2327 = in[2]? r2_4654 : r2_4653;
wire r3_2328;
assign r3_2328 = in[2]? r2_4656 : r2_4655;
wire r3_2329;
assign r3_2329 = in[2]? r2_4658 : r2_4657;
wire r3_2330;
assign r3_2330 = in[2]? r2_4660 : r2_4659;
wire r3_2331;
assign r3_2331 = in[2]? r2_4662 : r2_4661;
wire r3_2332;
assign r3_2332 = in[2]? r2_4664 : r2_4663;
wire r3_2333;
assign r3_2333 = in[2]? r2_4666 : r2_4665;
wire r3_2334;
assign r3_2334 = in[2]? r2_4668 : r2_4667;
wire r3_2335;
assign r3_2335 = in[2]? r2_4670 : r2_4669;
wire r3_2336;
assign r3_2336 = in[2]? r2_4672 : r2_4671;
wire r3_2337;
assign r3_2337 = in[2]? r2_4674 : r2_4673;
wire r3_2338;
assign r3_2338 = in[2]? r2_4676 : r2_4675;
wire r3_2339;
assign r3_2339 = in[2]? r2_4678 : r2_4677;
wire r3_2340;
assign r3_2340 = in[2]? r2_4680 : r2_4679;
wire r3_2341;
assign r3_2341 = in[2]? r2_4682 : r2_4681;
wire r3_2342;
assign r3_2342 = in[2]? r2_4684 : r2_4683;
wire r3_2343;
assign r3_2343 = in[2]? r2_4686 : r2_4685;
wire r3_2344;
assign r3_2344 = in[2]? r2_4688 : r2_4687;
wire r3_2345;
assign r3_2345 = in[2]? r2_4690 : r2_4689;
wire r3_2346;
assign r3_2346 = in[2]? r2_4692 : r2_4691;
wire r3_2347;
assign r3_2347 = in[2]? r2_4694 : r2_4693;
wire r3_2348;
assign r3_2348 = in[2]? r2_4696 : r2_4695;
wire r3_2349;
assign r3_2349 = in[2]? r2_4698 : r2_4697;
wire r3_2350;
assign r3_2350 = in[2]? r2_4700 : r2_4699;
wire r3_2351;
assign r3_2351 = in[2]? r2_4702 : r2_4701;
wire r3_2352;
assign r3_2352 = in[2]? r2_4704 : r2_4703;
wire r3_2353;
assign r3_2353 = in[2]? r2_4706 : r2_4705;
wire r3_2354;
assign r3_2354 = in[2]? r2_4708 : r2_4707;
wire r3_2355;
assign r3_2355 = in[2]? r2_4710 : r2_4709;
wire r3_2356;
assign r3_2356 = in[2]? r2_4712 : r2_4711;
wire r3_2357;
assign r3_2357 = in[2]? r2_4714 : r2_4713;
wire r3_2358;
assign r3_2358 = in[2]? r2_4716 : r2_4715;
wire r3_2359;
assign r3_2359 = in[2]? r2_4718 : r2_4717;
wire r3_2360;
assign r3_2360 = in[2]? r2_4720 : r2_4719;
wire r3_2361;
assign r3_2361 = in[2]? r2_4722 : r2_4721;
wire r3_2362;
assign r3_2362 = in[2]? r2_4724 : r2_4723;
wire r3_2363;
assign r3_2363 = in[2]? r2_4726 : r2_4725;
wire r3_2364;
assign r3_2364 = in[2]? r2_4728 : r2_4727;
wire r3_2365;
assign r3_2365 = in[2]? r2_4730 : r2_4729;
wire r3_2366;
assign r3_2366 = in[2]? r2_4732 : r2_4731;
wire r3_2367;
assign r3_2367 = in[2]? r2_4734 : r2_4733;
wire r3_2368;
assign r3_2368 = in[2]? r2_4736 : r2_4735;
wire r3_2369;
assign r3_2369 = in[2]? r2_4738 : r2_4737;
wire r3_2370;
assign r3_2370 = in[2]? r2_4740 : r2_4739;
wire r3_2371;
assign r3_2371 = in[2]? r2_4742 : r2_4741;
wire r3_2372;
assign r3_2372 = in[2]? r2_4744 : r2_4743;
wire r3_2373;
assign r3_2373 = in[2]? r2_4746 : r2_4745;
wire r3_2374;
assign r3_2374 = in[2]? r2_4748 : r2_4747;
wire r3_2375;
assign r3_2375 = in[2]? r2_4750 : r2_4749;
wire r3_2376;
assign r3_2376 = in[2]? r2_4752 : r2_4751;
wire r3_2377;
assign r3_2377 = in[2]? r2_4754 : r2_4753;
wire r3_2378;
assign r3_2378 = in[2]? r2_4756 : r2_4755;
wire r3_2379;
assign r3_2379 = in[2]? r2_4758 : r2_4757;
wire r3_2380;
assign r3_2380 = in[2]? r2_4760 : r2_4759;
wire r3_2381;
assign r3_2381 = in[2]? r2_4762 : r2_4761;
wire r3_2382;
assign r3_2382 = in[2]? r2_4764 : r2_4763;
wire r3_2383;
assign r3_2383 = in[2]? r2_4766 : r2_4765;
wire r3_2384;
assign r3_2384 = in[2]? r2_4768 : r2_4767;
wire r3_2385;
assign r3_2385 = in[2]? r2_4770 : r2_4769;
wire r3_2386;
assign r3_2386 = in[2]? r2_4772 : r2_4771;
wire r3_2387;
assign r3_2387 = in[2]? r2_4774 : r2_4773;
wire r3_2388;
assign r3_2388 = in[2]? r2_4776 : r2_4775;
wire r3_2389;
assign r3_2389 = in[2]? r2_4778 : r2_4777;
wire r3_2390;
assign r3_2390 = in[2]? r2_4780 : r2_4779;
wire r3_2391;
assign r3_2391 = in[2]? r2_4782 : r2_4781;
wire r3_2392;
assign r3_2392 = in[2]? r2_4784 : r2_4783;
wire r3_2393;
assign r3_2393 = in[2]? r2_4786 : r2_4785;
wire r3_2394;
assign r3_2394 = in[2]? r2_4788 : r2_4787;
wire r3_2395;
assign r3_2395 = in[2]? r2_4790 : r2_4789;
wire r3_2396;
assign r3_2396 = in[2]? r2_4792 : r2_4791;
wire r3_2397;
assign r3_2397 = in[2]? r2_4794 : r2_4793;
wire r3_2398;
assign r3_2398 = in[2]? r2_4796 : r2_4795;
wire r3_2399;
assign r3_2399 = in[2]? r2_4798 : r2_4797;
wire r3_2400;
assign r3_2400 = in[2]? r2_4800 : r2_4799;
wire r3_2401;
assign r3_2401 = in[2]? r2_4802 : r2_4801;
wire r3_2402;
assign r3_2402 = in[2]? r2_4804 : r2_4803;
wire r3_2403;
assign r3_2403 = in[2]? r2_4806 : r2_4805;
wire r3_2404;
assign r3_2404 = in[2]? r2_4808 : r2_4807;
wire r3_2405;
assign r3_2405 = in[2]? r2_4810 : r2_4809;
wire r3_2406;
assign r3_2406 = in[2]? r2_4812 : r2_4811;
wire r3_2407;
assign r3_2407 = in[2]? r2_4814 : r2_4813;
wire r3_2408;
assign r3_2408 = in[2]? r2_4816 : r2_4815;
wire r3_2409;
assign r3_2409 = in[2]? r2_4818 : r2_4817;
wire r3_2410;
assign r3_2410 = in[2]? r2_4820 : r2_4819;
wire r3_2411;
assign r3_2411 = in[2]? r2_4822 : r2_4821;
wire r3_2412;
assign r3_2412 = in[2]? r2_4824 : r2_4823;
wire r3_2413;
assign r3_2413 = in[2]? r2_4826 : r2_4825;
wire r3_2414;
assign r3_2414 = in[2]? r2_4828 : r2_4827;
wire r3_2415;
assign r3_2415 = in[2]? r2_4830 : r2_4829;
wire r3_2416;
assign r3_2416 = in[2]? r2_4832 : r2_4831;
wire r3_2417;
assign r3_2417 = in[2]? r2_4834 : r2_4833;
wire r3_2418;
assign r3_2418 = in[2]? r2_4836 : r2_4835;
wire r3_2419;
assign r3_2419 = in[2]? r2_4838 : r2_4837;
wire r3_2420;
assign r3_2420 = in[2]? r2_4840 : r2_4839;
wire r3_2421;
assign r3_2421 = in[2]? r2_4842 : r2_4841;
wire r3_2422;
assign r3_2422 = in[2]? r2_4844 : r2_4843;
wire r3_2423;
assign r3_2423 = in[2]? r2_4846 : r2_4845;
wire r3_2424;
assign r3_2424 = in[2]? r2_4848 : r2_4847;
wire r3_2425;
assign r3_2425 = in[2]? r2_4850 : r2_4849;
wire r3_2426;
assign r3_2426 = in[2]? r2_4852 : r2_4851;
wire r3_2427;
assign r3_2427 = in[2]? r2_4854 : r2_4853;
wire r3_2428;
assign r3_2428 = in[2]? r2_4856 : r2_4855;
wire r3_2429;
assign r3_2429 = in[2]? r2_4858 : r2_4857;
wire r3_2430;
assign r3_2430 = in[2]? r2_4860 : r2_4859;
wire r3_2431;
assign r3_2431 = in[2]? r2_4862 : r2_4861;
wire r3_2432;
assign r3_2432 = in[2]? r2_4864 : r2_4863;
wire r3_2433;
assign r3_2433 = in[2]? r2_4866 : r2_4865;
wire r3_2434;
assign r3_2434 = in[2]? r2_4868 : r2_4867;
wire r3_2435;
assign r3_2435 = in[2]? r2_4870 : r2_4869;
wire r3_2436;
assign r3_2436 = in[2]? r2_4872 : r2_4871;
wire r3_2437;
assign r3_2437 = in[2]? r2_4874 : r2_4873;
wire r3_2438;
assign r3_2438 = in[2]? r2_4876 : r2_4875;
wire r3_2439;
assign r3_2439 = in[2]? r2_4878 : r2_4877;
wire r3_2440;
assign r3_2440 = in[2]? r2_4880 : r2_4879;
wire r3_2441;
assign r3_2441 = in[2]? r2_4882 : r2_4881;
wire r3_2442;
assign r3_2442 = in[2]? r2_4884 : r2_4883;
wire r3_2443;
assign r3_2443 = in[2]? r2_4886 : r2_4885;
wire r3_2444;
assign r3_2444 = in[2]? r2_4888 : r2_4887;
wire r3_2445;
assign r3_2445 = in[2]? r2_4890 : r2_4889;
wire r3_2446;
assign r3_2446 = in[2]? r2_4892 : r2_4891;
wire r3_2447;
assign r3_2447 = in[2]? r2_4894 : r2_4893;
wire r3_2448;
assign r3_2448 = in[2]? r2_4896 : r2_4895;
wire r3_2449;
assign r3_2449 = in[2]? r2_4898 : r2_4897;
wire r3_2450;
assign r3_2450 = in[2]? r2_4900 : r2_4899;
wire r3_2451;
assign r3_2451 = in[2]? r2_4902 : r2_4901;
wire r3_2452;
assign r3_2452 = in[2]? r2_4904 : r2_4903;
wire r3_2453;
assign r3_2453 = in[2]? r2_4906 : r2_4905;
wire r3_2454;
assign r3_2454 = in[2]? r2_4908 : r2_4907;
wire r3_2455;
assign r3_2455 = in[2]? r2_4910 : r2_4909;
wire r3_2456;
assign r3_2456 = in[2]? r2_4912 : r2_4911;
wire r3_2457;
assign r3_2457 = in[2]? r2_4914 : r2_4913;
wire r3_2458;
assign r3_2458 = in[2]? r2_4916 : r2_4915;
wire r3_2459;
assign r3_2459 = in[2]? r2_4918 : r2_4917;
wire r3_2460;
assign r3_2460 = in[2]? r2_4920 : r2_4919;
wire r3_2461;
assign r3_2461 = in[2]? r2_4922 : r2_4921;
wire r3_2462;
assign r3_2462 = in[2]? r2_4924 : r2_4923;
wire r3_2463;
assign r3_2463 = in[2]? r2_4926 : r2_4925;
wire r3_2464;
assign r3_2464 = in[2]? r2_4928 : r2_4927;
wire r3_2465;
assign r3_2465 = in[2]? r2_4930 : r2_4929;
wire r3_2466;
assign r3_2466 = in[2]? r2_4932 : r2_4931;
wire r3_2467;
assign r3_2467 = in[2]? r2_4934 : r2_4933;
wire r3_2468;
assign r3_2468 = in[2]? r2_4936 : r2_4935;
wire r3_2469;
assign r3_2469 = in[2]? r2_4938 : r2_4937;
wire r3_2470;
assign r3_2470 = in[2]? r2_4940 : r2_4939;
wire r3_2471;
assign r3_2471 = in[2]? r2_4942 : r2_4941;
wire r3_2472;
assign r3_2472 = in[2]? r2_4944 : r2_4943;
wire r3_2473;
assign r3_2473 = in[2]? r2_4946 : r2_4945;
wire r3_2474;
assign r3_2474 = in[2]? r2_4948 : r2_4947;
wire r3_2475;
assign r3_2475 = in[2]? r2_4950 : r2_4949;
wire r3_2476;
assign r3_2476 = in[2]? r2_4952 : r2_4951;
wire r3_2477;
assign r3_2477 = in[2]? r2_4954 : r2_4953;
wire r3_2478;
assign r3_2478 = in[2]? r2_4956 : r2_4955;
wire r3_2479;
assign r3_2479 = in[2]? r2_4958 : r2_4957;
wire r3_2480;
assign r3_2480 = in[2]? r2_4960 : r2_4959;
wire r3_2481;
assign r3_2481 = in[2]? r2_4962 : r2_4961;
wire r3_2482;
assign r3_2482 = in[2]? r2_4964 : r2_4963;
wire r3_2483;
assign r3_2483 = in[2]? r2_4966 : r2_4965;
wire r3_2484;
assign r3_2484 = in[2]? r2_4968 : r2_4967;
wire r3_2485;
assign r3_2485 = in[2]? r2_4970 : r2_4969;
wire r3_2486;
assign r3_2486 = in[2]? r2_4972 : r2_4971;
wire r3_2487;
assign r3_2487 = in[2]? r2_4974 : r2_4973;
wire r3_2488;
assign r3_2488 = in[2]? r2_4976 : r2_4975;
wire r3_2489;
assign r3_2489 = in[2]? r2_4978 : r2_4977;
wire r3_2490;
assign r3_2490 = in[2]? r2_4980 : r2_4979;
wire r3_2491;
assign r3_2491 = in[2]? r2_4982 : r2_4981;
wire r3_2492;
assign r3_2492 = in[2]? r2_4984 : r2_4983;
wire r3_2493;
assign r3_2493 = in[2]? r2_4986 : r2_4985;
wire r3_2494;
assign r3_2494 = in[2]? r2_4988 : r2_4987;
wire r3_2495;
assign r3_2495 = in[2]? r2_4990 : r2_4989;
wire r3_2496;
assign r3_2496 = in[2]? r2_4992 : r2_4991;
wire r3_2497;
assign r3_2497 = in[2]? r2_4994 : r2_4993;
wire r3_2498;
assign r3_2498 = in[2]? r2_4996 : r2_4995;
wire r3_2499;
assign r3_2499 = in[2]? r2_4998 : r2_4997;
wire r3_2500;
assign r3_2500 = in[2]? r2_5000 : r2_4999;
wire r3_2501;
assign r3_2501 = in[2]? r2_5002 : r2_5001;
wire r3_2502;
assign r3_2502 = in[2]? r2_5004 : r2_5003;
wire r3_2503;
assign r3_2503 = in[2]? r2_5006 : r2_5005;
wire r3_2504;
assign r3_2504 = in[2]? r2_5008 : r2_5007;
wire r3_2505;
assign r3_2505 = in[2]? r2_5010 : r2_5009;
wire r3_2506;
assign r3_2506 = in[2]? r2_5012 : r2_5011;
wire r3_2507;
assign r3_2507 = in[2]? r2_5014 : r2_5013;
wire r3_2508;
assign r3_2508 = in[2]? r2_5016 : r2_5015;
wire r3_2509;
assign r3_2509 = in[2]? r2_5018 : r2_5017;
wire r3_2510;
assign r3_2510 = in[2]? r2_5020 : r2_5019;
wire r3_2511;
assign r3_2511 = in[2]? r2_5022 : r2_5021;
wire r3_2512;
assign r3_2512 = in[2]? r2_5024 : r2_5023;
wire r3_2513;
assign r3_2513 = in[2]? r2_5026 : r2_5025;
wire r3_2514;
assign r3_2514 = in[2]? r2_5028 : r2_5027;
wire r3_2515;
assign r3_2515 = in[2]? r2_5030 : r2_5029;
wire r3_2516;
assign r3_2516 = in[2]? r2_5032 : r2_5031;
wire r3_2517;
assign r3_2517 = in[2]? r2_5034 : r2_5033;
wire r3_2518;
assign r3_2518 = in[2]? r2_5036 : r2_5035;
wire r3_2519;
assign r3_2519 = in[2]? r2_5038 : r2_5037;
wire r3_2520;
assign r3_2520 = in[2]? r2_5040 : r2_5039;
wire r3_2521;
assign r3_2521 = in[2]? r2_5042 : r2_5041;
wire r3_2522;
assign r3_2522 = in[2]? r2_5044 : r2_5043;
wire r3_2523;
assign r3_2523 = in[2]? r2_5046 : r2_5045;
wire r3_2524;
assign r3_2524 = in[2]? r2_5048 : r2_5047;
wire r3_2525;
assign r3_2525 = in[2]? r2_5050 : r2_5049;
wire r3_2526;
assign r3_2526 = in[2]? r2_5052 : r2_5051;
wire r3_2527;
assign r3_2527 = in[2]? r2_5054 : r2_5053;
wire r3_2528;
assign r3_2528 = in[2]? r2_5056 : r2_5055;
wire r3_2529;
assign r3_2529 = in[2]? r2_5058 : r2_5057;
wire r3_2530;
assign r3_2530 = in[2]? r2_5060 : r2_5059;
wire r3_2531;
assign r3_2531 = in[2]? r2_5062 : r2_5061;
wire r3_2532;
assign r3_2532 = in[2]? r2_5064 : r2_5063;
wire r3_2533;
assign r3_2533 = in[2]? r2_5066 : r2_5065;
wire r3_2534;
assign r3_2534 = in[2]? r2_5068 : r2_5067;
wire r3_2535;
assign r3_2535 = in[2]? r2_5070 : r2_5069;
wire r3_2536;
assign r3_2536 = in[2]? r2_5072 : r2_5071;
wire r3_2537;
assign r3_2537 = in[2]? r2_5074 : r2_5073;
wire r3_2538;
assign r3_2538 = in[2]? r2_5076 : r2_5075;
wire r3_2539;
assign r3_2539 = in[2]? r2_5078 : r2_5077;
wire r3_2540;
assign r3_2540 = in[2]? r2_5080 : r2_5079;
wire r3_2541;
assign r3_2541 = in[2]? r2_5082 : r2_5081;
wire r3_2542;
assign r3_2542 = in[2]? r2_5084 : r2_5083;
wire r3_2543;
assign r3_2543 = in[2]? r2_5086 : r2_5085;
wire r3_2544;
assign r3_2544 = in[2]? r2_5088 : r2_5087;
wire r3_2545;
assign r3_2545 = in[2]? r2_5090 : r2_5089;
wire r3_2546;
assign r3_2546 = in[2]? r2_5092 : r2_5091;
wire r3_2547;
assign r3_2547 = in[2]? r2_5094 : r2_5093;
wire r3_2548;
assign r3_2548 = in[2]? r2_5096 : r2_5095;
wire r3_2549;
assign r3_2549 = in[2]? r2_5098 : r2_5097;
wire r3_2550;
assign r3_2550 = in[2]? r2_5100 : r2_5099;
wire r3_2551;
assign r3_2551 = in[2]? r2_5102 : r2_5101;
wire r3_2552;
assign r3_2552 = in[2]? r2_5104 : r2_5103;
wire r3_2553;
assign r3_2553 = in[2]? r2_5106 : r2_5105;
wire r3_2554;
assign r3_2554 = in[2]? r2_5108 : r2_5107;
wire r3_2555;
assign r3_2555 = in[2]? r2_5110 : r2_5109;
wire r3_2556;
assign r3_2556 = in[2]? r2_5112 : r2_5111;
wire r3_2557;
assign r3_2557 = in[2]? r2_5114 : r2_5113;
wire r3_2558;
assign r3_2558 = in[2]? r2_5116 : r2_5115;
wire r3_2559;
assign r3_2559 = in[2]? r2_5118 : r2_5117;
wire r3_2560;
assign r3_2560 = in[2]? r2_5120 : r2_5119;
wire r3_2561;
assign r3_2561 = in[2]? r2_5122 : r2_5121;
wire r3_2562;
assign r3_2562 = in[2]? r2_5124 : r2_5123;
wire r3_2563;
assign r3_2563 = in[2]? r2_5126 : r2_5125;
wire r3_2564;
assign r3_2564 = in[2]? r2_5128 : r2_5127;
wire r3_2565;
assign r3_2565 = in[2]? r2_5130 : r2_5129;
wire r3_2566;
assign r3_2566 = in[2]? r2_5132 : r2_5131;
wire r3_2567;
assign r3_2567 = in[2]? r2_5134 : r2_5133;
wire r3_2568;
assign r3_2568 = in[2]? r2_5136 : r2_5135;
wire r4_1;
assign r4_1 = in[3]? r3_2 : r3_1;
wire r4_2;
assign r4_2 = in[3]? r3_4 : r3_3;
wire r4_3;
assign r4_3 = in[3]? r3_6 : r3_5;
wire r4_4;
assign r4_4 = in[3]? r3_8 : r3_7;
wire r4_5;
assign r4_5 = in[3]? r3_10 : r3_9;
wire r4_6;
assign r4_6 = in[3]? r3_12 : r3_11;
wire r4_7;
assign r4_7 = in[3]? r3_14 : r3_13;
wire r4_8;
assign r4_8 = in[3]? r3_16 : r3_15;
wire r4_9;
assign r4_9 = in[3]? r3_18 : r3_17;
wire r4_10;
assign r4_10 = in[3]? r3_20 : r3_19;
wire r4_11;
assign r4_11 = in[3]? r3_22 : r3_21;
wire r4_12;
assign r4_12 = in[3]? r3_24 : r3_23;
wire r4_13;
assign r4_13 = in[3]? r3_26 : r3_25;
wire r4_14;
assign r4_14 = in[3]? r3_28 : r3_27;
wire r4_15;
assign r4_15 = in[3]? r3_30 : r3_29;
wire r4_16;
assign r4_16 = in[3]? r3_32 : r3_31;
wire r4_17;
assign r4_17 = in[3]? r3_34 : r3_33;
wire r4_18;
assign r4_18 = in[3]? r3_36 : r3_35;
wire r4_19;
assign r4_19 = in[3]? r3_38 : r3_37;
wire r4_20;
assign r4_20 = in[3]? r3_40 : r3_39;
wire r4_21;
assign r4_21 = in[3]? r3_42 : r3_41;
wire r4_22;
assign r4_22 = in[3]? r3_44 : r3_43;
wire r4_23;
assign r4_23 = in[3]? r3_46 : r3_45;
wire r4_24;
assign r4_24 = in[3]? r3_48 : r3_47;
wire r4_25;
assign r4_25 = in[3]? r3_50 : r3_49;
wire r4_26;
assign r4_26 = in[3]? r3_52 : r3_51;
wire r4_27;
assign r4_27 = in[3]? r3_54 : r3_53;
wire r4_28;
assign r4_28 = in[3]? r3_56 : r3_55;
wire r4_29;
assign r4_29 = in[3]? r3_58 : r3_57;
wire r4_30;
assign r4_30 = in[3]? r3_60 : r3_59;
wire r4_31;
assign r4_31 = in[3]? r3_62 : r3_61;
wire r4_32;
assign r4_32 = in[3]? r3_64 : r3_63;
wire r4_33;
assign r4_33 = in[3]? r3_66 : r3_65;
wire r4_34;
assign r4_34 = in[3]? r3_68 : r3_67;
wire r4_35;
assign r4_35 = in[3]? r3_70 : r3_69;
wire r4_36;
assign r4_36 = in[3]? r3_72 : r3_71;
wire r4_37;
assign r4_37 = in[3]? r3_74 : r3_73;
wire r4_38;
assign r4_38 = in[3]? r3_76 : r3_75;
wire r4_39;
assign r4_39 = in[3]? r3_78 : r3_77;
wire r4_40;
assign r4_40 = in[3]? r3_80 : r3_79;
wire r4_41;
assign r4_41 = in[3]? r3_82 : r3_81;
wire r4_42;
assign r4_42 = in[3]? r3_84 : r3_83;
wire r4_43;
assign r4_43 = in[3]? r3_86 : r3_85;
wire r4_44;
assign r4_44 = in[3]? r3_88 : r3_87;
wire r4_45;
assign r4_45 = in[3]? r3_90 : r3_89;
wire r4_46;
assign r4_46 = in[3]? r3_92 : r3_91;
wire r4_47;
assign r4_47 = in[3]? r3_94 : r3_93;
wire r4_48;
assign r4_48 = in[3]? r3_96 : r3_95;
wire r4_49;
assign r4_49 = in[3]? r3_98 : r3_97;
wire r4_50;
assign r4_50 = in[3]? r3_100 : r3_99;
wire r4_51;
assign r4_51 = in[3]? r3_102 : r3_101;
wire r4_52;
assign r4_52 = in[3]? r3_104 : r3_103;
wire r4_53;
assign r4_53 = in[3]? r3_106 : r3_105;
wire r4_54;
assign r4_54 = in[3]? r3_108 : r3_107;
wire r4_55;
assign r4_55 = in[3]? r3_110 : r3_109;
wire r4_56;
assign r4_56 = in[3]? r3_112 : r3_111;
wire r4_57;
assign r4_57 = in[3]? r3_114 : r3_113;
wire r4_58;
assign r4_58 = in[3]? r3_116 : r3_115;
wire r4_59;
assign r4_59 = in[3]? r3_118 : r3_117;
wire r4_60;
assign r4_60 = in[3]? r3_120 : r3_119;
wire r4_61;
assign r4_61 = in[3]? r3_122 : r3_121;
wire r4_62;
assign r4_62 = in[3]? r3_124 : r3_123;
wire r4_63;
assign r4_63 = in[3]? r3_126 : r3_125;
wire r4_64;
assign r4_64 = in[3]? r3_128 : r3_127;
wire r4_65;
assign r4_65 = in[3]? r3_130 : r3_129;
wire r4_66;
assign r4_66 = in[3]? r3_132 : r3_131;
wire r4_67;
assign r4_67 = in[3]? r3_134 : r3_133;
wire r4_68;
assign r4_68 = in[3]? r3_136 : r3_135;
wire r4_69;
assign r4_69 = in[3]? r3_138 : r3_137;
wire r4_70;
assign r4_70 = in[3]? r3_140 : r3_139;
wire r4_71;
assign r4_71 = in[3]? r3_142 : r3_141;
wire r4_72;
assign r4_72 = in[3]? r3_144 : r3_143;
wire r4_73;
assign r4_73 = in[3]? r3_146 : r3_145;
wire r4_74;
assign r4_74 = in[3]? r3_148 : r3_147;
wire r4_75;
assign r4_75 = in[3]? r3_150 : r3_149;
wire r4_76;
assign r4_76 = in[3]? r3_152 : r3_151;
wire r4_77;
assign r4_77 = in[3]? r3_154 : r3_153;
wire r4_78;
assign r4_78 = in[3]? r3_156 : r3_155;
wire r4_79;
assign r4_79 = in[3]? r3_158 : r3_157;
wire r4_80;
assign r4_80 = in[3]? r3_160 : r3_159;
wire r4_81;
assign r4_81 = in[3]? r3_162 : r3_161;
wire r4_82;
assign r4_82 = in[3]? r3_164 : r3_163;
wire r4_83;
assign r4_83 = in[3]? r3_166 : r3_165;
wire r4_84;
assign r4_84 = in[3]? r3_168 : r3_167;
wire r4_85;
assign r4_85 = in[3]? r3_170 : r3_169;
wire r4_86;
assign r4_86 = in[3]? r3_172 : r3_171;
wire r4_87;
assign r4_87 = in[3]? r3_174 : r3_173;
wire r4_88;
assign r4_88 = in[3]? r3_176 : r3_175;
wire r4_89;
assign r4_89 = in[3]? r3_178 : r3_177;
wire r4_90;
assign r4_90 = in[3]? r3_180 : r3_179;
wire r4_91;
assign r4_91 = in[3]? r3_182 : r3_181;
wire r4_92;
assign r4_92 = in[3]? r3_184 : r3_183;
wire r4_93;
assign r4_93 = in[3]? r3_186 : r3_185;
wire r4_94;
assign r4_94 = in[3]? r3_188 : r3_187;
wire r4_95;
assign r4_95 = in[3]? r3_190 : r3_189;
wire r4_96;
assign r4_96 = in[3]? r3_192 : r3_191;
wire r4_97;
assign r4_97 = in[3]? r3_194 : r3_193;
wire r4_98;
assign r4_98 = in[3]? r3_196 : r3_195;
wire r4_99;
assign r4_99 = in[3]? r3_198 : r3_197;
wire r4_100;
assign r4_100 = in[3]? r3_200 : r3_199;
wire r4_101;
assign r4_101 = in[3]? r3_202 : r3_201;
wire r4_102;
assign r4_102 = in[3]? r3_204 : r3_203;
wire r4_103;
assign r4_103 = in[3]? r3_206 : r3_205;
wire r4_104;
assign r4_104 = in[3]? r3_208 : r3_207;
wire r4_105;
assign r4_105 = in[3]? r3_210 : r3_209;
wire r4_106;
assign r4_106 = in[3]? r3_212 : r3_211;
wire r4_107;
assign r4_107 = in[3]? r3_214 : r3_213;
wire r4_108;
assign r4_108 = in[3]? r3_216 : r3_215;
wire r4_109;
assign r4_109 = in[3]? r3_218 : r3_217;
wire r4_110;
assign r4_110 = in[3]? r3_220 : r3_219;
wire r4_111;
assign r4_111 = in[3]? r3_222 : r3_221;
wire r4_112;
assign r4_112 = in[3]? r3_224 : r3_223;
wire r4_113;
assign r4_113 = in[3]? r3_226 : r3_225;
wire r4_114;
assign r4_114 = in[3]? r3_228 : r3_227;
wire r4_115;
assign r4_115 = in[3]? r3_230 : r3_229;
wire r4_116;
assign r4_116 = in[3]? r3_232 : r3_231;
wire r4_117;
assign r4_117 = in[3]? r3_234 : r3_233;
wire r4_118;
assign r4_118 = in[3]? r3_236 : r3_235;
wire r4_119;
assign r4_119 = in[3]? r3_238 : r3_237;
wire r4_120;
assign r4_120 = in[3]? r3_240 : r3_239;
wire r4_121;
assign r4_121 = in[3]? r3_242 : r3_241;
wire r4_122;
assign r4_122 = in[3]? r3_244 : r3_243;
wire r4_123;
assign r4_123 = in[3]? r3_246 : r3_245;
wire r4_124;
assign r4_124 = in[3]? r3_248 : r3_247;
wire r4_125;
assign r4_125 = in[3]? r3_250 : r3_249;
wire r4_126;
assign r4_126 = in[3]? r3_252 : r3_251;
wire r4_127;
assign r4_127 = in[3]? r3_254 : r3_253;
wire r4_128;
assign r4_128 = in[3]? r3_256 : r3_255;
wire r4_129;
assign r4_129 = in[3]? r3_258 : r3_257;
wire r4_130;
assign r4_130 = in[3]? r3_260 : r3_259;
wire r4_131;
assign r4_131 = in[3]? r3_262 : r3_261;
wire r4_132;
assign r4_132 = in[3]? r3_264 : r3_263;
wire r4_133;
assign r4_133 = in[3]? r3_266 : r3_265;
wire r4_134;
assign r4_134 = in[3]? r3_268 : r3_267;
wire r4_135;
assign r4_135 = in[3]? r3_270 : r3_269;
wire r4_136;
assign r4_136 = in[3]? r3_272 : r3_271;
wire r4_137;
assign r4_137 = in[3]? r3_274 : r3_273;
wire r4_138;
assign r4_138 = in[3]? r3_276 : r3_275;
wire r4_139;
assign r4_139 = in[3]? r3_278 : r3_277;
wire r4_140;
assign r4_140 = in[3]? r3_280 : r3_279;
wire r4_141;
assign r4_141 = in[3]? r3_282 : r3_281;
wire r4_142;
assign r4_142 = in[3]? r3_284 : r3_283;
wire r4_143;
assign r4_143 = in[3]? r3_286 : r3_285;
wire r4_144;
assign r4_144 = in[3]? r3_288 : r3_287;
wire r4_145;
assign r4_145 = in[3]? r3_290 : r3_289;
wire r4_146;
assign r4_146 = in[3]? r3_292 : r3_291;
wire r4_147;
assign r4_147 = in[3]? r3_294 : r3_293;
wire r4_148;
assign r4_148 = in[3]? r3_296 : r3_295;
wire r4_149;
assign r4_149 = in[3]? r3_298 : r3_297;
wire r4_150;
assign r4_150 = in[3]? r3_300 : r3_299;
wire r4_151;
assign r4_151 = in[3]? r3_302 : r3_301;
wire r4_152;
assign r4_152 = in[3]? r3_304 : r3_303;
wire r4_153;
assign r4_153 = in[3]? r3_306 : r3_305;
wire r4_154;
assign r4_154 = in[3]? r3_308 : r3_307;
wire r4_155;
assign r4_155 = in[3]? r3_310 : r3_309;
wire r4_156;
assign r4_156 = in[3]? r3_312 : r3_311;
wire r4_157;
assign r4_157 = in[3]? r3_314 : r3_313;
wire r4_158;
assign r4_158 = in[3]? r3_316 : r3_315;
wire r4_159;
assign r4_159 = in[3]? r3_318 : r3_317;
wire r4_160;
assign r4_160 = in[3]? r3_320 : r3_319;
wire r4_161;
assign r4_161 = in[3]? r3_322 : r3_321;
wire r4_162;
assign r4_162 = in[3]? r3_324 : r3_323;
wire r4_163;
assign r4_163 = in[3]? r3_326 : r3_325;
wire r4_164;
assign r4_164 = in[3]? r3_328 : r3_327;
wire r4_165;
assign r4_165 = in[3]? r3_330 : r3_329;
wire r4_166;
assign r4_166 = in[3]? r3_332 : r3_331;
wire r4_167;
assign r4_167 = in[3]? r3_334 : r3_333;
wire r4_168;
assign r4_168 = in[3]? r3_336 : r3_335;
wire r4_169;
assign r4_169 = in[3]? r3_338 : r3_337;
wire r4_170;
assign r4_170 = in[3]? r3_340 : r3_339;
wire r4_171;
assign r4_171 = in[3]? r3_342 : r3_341;
wire r4_172;
assign r4_172 = in[3]? r3_344 : r3_343;
wire r4_173;
assign r4_173 = in[3]? r3_346 : r3_345;
wire r4_174;
assign r4_174 = in[3]? r3_348 : r3_347;
wire r4_175;
assign r4_175 = in[3]? r3_350 : r3_349;
wire r4_176;
assign r4_176 = in[3]? r3_352 : r3_351;
wire r4_177;
assign r4_177 = in[3]? r3_354 : r3_353;
wire r4_178;
assign r4_178 = in[3]? r3_356 : r3_355;
wire r4_179;
assign r4_179 = in[3]? r3_358 : r3_357;
wire r4_180;
assign r4_180 = in[3]? r3_360 : r3_359;
wire r4_181;
assign r4_181 = in[3]? r3_362 : r3_361;
wire r4_182;
assign r4_182 = in[3]? r3_364 : r3_363;
wire r4_183;
assign r4_183 = in[3]? r3_366 : r3_365;
wire r4_184;
assign r4_184 = in[3]? r3_368 : r3_367;
wire r4_185;
assign r4_185 = in[3]? r3_370 : r3_369;
wire r4_186;
assign r4_186 = in[3]? r3_372 : r3_371;
wire r4_187;
assign r4_187 = in[3]? r3_374 : r3_373;
wire r4_188;
assign r4_188 = in[3]? r3_376 : r3_375;
wire r4_189;
assign r4_189 = in[3]? r3_378 : r3_377;
wire r4_190;
assign r4_190 = in[3]? r3_380 : r3_379;
wire r4_191;
assign r4_191 = in[3]? r3_382 : r3_381;
wire r4_192;
assign r4_192 = in[3]? r3_384 : r3_383;
wire r4_193;
assign r4_193 = in[3]? r3_386 : r3_385;
wire r4_194;
assign r4_194 = in[3]? r3_388 : r3_387;
wire r4_195;
assign r4_195 = in[3]? r3_390 : r3_389;
wire r4_196;
assign r4_196 = in[3]? r3_392 : r3_391;
wire r4_197;
assign r4_197 = in[3]? r3_394 : r3_393;
wire r4_198;
assign r4_198 = in[3]? r3_396 : r3_395;
wire r4_199;
assign r4_199 = in[3]? r3_398 : r3_397;
wire r4_200;
assign r4_200 = in[3]? r3_400 : r3_399;
wire r4_201;
assign r4_201 = in[3]? r3_402 : r3_401;
wire r4_202;
assign r4_202 = in[3]? r3_404 : r3_403;
wire r4_203;
assign r4_203 = in[3]? r3_406 : r3_405;
wire r4_204;
assign r4_204 = in[3]? r3_408 : r3_407;
wire r4_205;
assign r4_205 = in[3]? r3_410 : r3_409;
wire r4_206;
assign r4_206 = in[3]? r3_412 : r3_411;
wire r4_207;
assign r4_207 = in[3]? r3_414 : r3_413;
wire r4_208;
assign r4_208 = in[3]? r3_416 : r3_415;
wire r4_209;
assign r4_209 = in[3]? r3_418 : r3_417;
wire r4_210;
assign r4_210 = in[3]? r3_420 : r3_419;
wire r4_211;
assign r4_211 = in[3]? r3_422 : r3_421;
wire r4_212;
assign r4_212 = in[3]? r3_424 : r3_423;
wire r4_213;
assign r4_213 = in[3]? r3_426 : r3_425;
wire r4_214;
assign r4_214 = in[3]? r3_428 : r3_427;
wire r4_215;
assign r4_215 = in[3]? r3_430 : r3_429;
wire r4_216;
assign r4_216 = in[3]? r3_432 : r3_431;
wire r4_217;
assign r4_217 = in[3]? r3_434 : r3_433;
wire r4_218;
assign r4_218 = in[3]? r3_436 : r3_435;
wire r4_219;
assign r4_219 = in[3]? r3_438 : r3_437;
wire r4_220;
assign r4_220 = in[3]? r3_440 : r3_439;
wire r4_221;
assign r4_221 = in[3]? r3_442 : r3_441;
wire r4_222;
assign r4_222 = in[3]? r3_444 : r3_443;
wire r4_223;
assign r4_223 = in[3]? r3_446 : r3_445;
wire r4_224;
assign r4_224 = in[3]? r3_448 : r3_447;
wire r4_225;
assign r4_225 = in[3]? r3_450 : r3_449;
wire r4_226;
assign r4_226 = in[3]? r3_452 : r3_451;
wire r4_227;
assign r4_227 = in[3]? r3_454 : r3_453;
wire r4_228;
assign r4_228 = in[3]? r3_456 : r3_455;
wire r4_229;
assign r4_229 = in[3]? r3_458 : r3_457;
wire r4_230;
assign r4_230 = in[3]? r3_460 : r3_459;
wire r4_231;
assign r4_231 = in[3]? r3_462 : r3_461;
wire r4_232;
assign r4_232 = in[3]? r3_464 : r3_463;
wire r4_233;
assign r4_233 = in[3]? r3_466 : r3_465;
wire r4_234;
assign r4_234 = in[3]? r3_468 : r3_467;
wire r4_235;
assign r4_235 = in[3]? r3_470 : r3_469;
wire r4_236;
assign r4_236 = in[3]? r3_472 : r3_471;
wire r4_237;
assign r4_237 = in[3]? r3_474 : r3_473;
wire r4_238;
assign r4_238 = in[3]? r3_476 : r3_475;
wire r4_239;
assign r4_239 = in[3]? r3_478 : r3_477;
wire r4_240;
assign r4_240 = in[3]? r3_480 : r3_479;
wire r4_241;
assign r4_241 = in[3]? r3_482 : r3_481;
wire r4_242;
assign r4_242 = in[3]? r3_484 : r3_483;
wire r4_243;
assign r4_243 = in[3]? r3_486 : r3_485;
wire r4_244;
assign r4_244 = in[3]? r3_488 : r3_487;
wire r4_245;
assign r4_245 = in[3]? r3_490 : r3_489;
wire r4_246;
assign r4_246 = in[3]? r3_492 : r3_491;
wire r4_247;
assign r4_247 = in[3]? r3_494 : r3_493;
wire r4_248;
assign r4_248 = in[3]? r3_496 : r3_495;
wire r4_249;
assign r4_249 = in[3]? r3_498 : r3_497;
wire r4_250;
assign r4_250 = in[3]? r3_500 : r3_499;
wire r4_251;
assign r4_251 = in[3]? r3_502 : r3_501;
wire r4_252;
assign r4_252 = in[3]? r3_504 : r3_503;
wire r4_253;
assign r4_253 = in[3]? r3_506 : r3_505;
wire r4_254;
assign r4_254 = in[3]? r3_508 : r3_507;
wire r4_255;
assign r4_255 = in[3]? r3_510 : r3_509;
wire r4_256;
assign r4_256 = in[3]? r3_512 : r3_511;
wire r4_257;
assign r4_257 = in[3]? r3_514 : r3_513;
wire r4_258;
assign r4_258 = in[3]? r3_516 : r3_515;
wire r4_259;
assign r4_259 = in[3]? r3_518 : r3_517;
wire r4_260;
assign r4_260 = in[3]? r3_520 : r3_519;
wire r4_261;
assign r4_261 = in[3]? r3_522 : r3_521;
wire r4_262;
assign r4_262 = in[3]? r3_524 : r3_523;
wire r4_263;
assign r4_263 = in[3]? r3_526 : r3_525;
wire r4_264;
assign r4_264 = in[3]? r3_528 : r3_527;
wire r4_265;
assign r4_265 = in[3]? r3_530 : r3_529;
wire r4_266;
assign r4_266 = in[3]? r3_532 : r3_531;
wire r4_267;
assign r4_267 = in[3]? r3_534 : r3_533;
wire r4_268;
assign r4_268 = in[3]? r3_536 : r3_535;
wire r4_269;
assign r4_269 = in[3]? r3_538 : r3_537;
wire r4_270;
assign r4_270 = in[3]? r3_540 : r3_539;
wire r4_271;
assign r4_271 = in[3]? r3_542 : r3_541;
wire r4_272;
assign r4_272 = in[3]? r3_544 : r3_543;
wire r4_273;
assign r4_273 = in[3]? r3_546 : r3_545;
wire r4_274;
assign r4_274 = in[3]? r3_548 : r3_547;
wire r4_275;
assign r4_275 = in[3]? r3_550 : r3_549;
wire r4_276;
assign r4_276 = in[3]? r3_552 : r3_551;
wire r4_277;
assign r4_277 = in[3]? r3_554 : r3_553;
wire r4_278;
assign r4_278 = in[3]? r3_556 : r3_555;
wire r4_279;
assign r4_279 = in[3]? r3_558 : r3_557;
wire r4_280;
assign r4_280 = in[3]? r3_560 : r3_559;
wire r4_281;
assign r4_281 = in[3]? r3_562 : r3_561;
wire r4_282;
assign r4_282 = in[3]? r3_564 : r3_563;
wire r4_283;
assign r4_283 = in[3]? r3_566 : r3_565;
wire r4_284;
assign r4_284 = in[3]? r3_568 : r3_567;
wire r4_285;
assign r4_285 = in[3]? r3_570 : r3_569;
wire r4_286;
assign r4_286 = in[3]? r3_572 : r3_571;
wire r4_287;
assign r4_287 = in[3]? r3_574 : r3_573;
wire r4_288;
assign r4_288 = in[3]? r3_576 : r3_575;
wire r4_289;
assign r4_289 = in[3]? r3_578 : r3_577;
wire r4_290;
assign r4_290 = in[3]? r3_580 : r3_579;
wire r4_291;
assign r4_291 = in[3]? r3_582 : r3_581;
wire r4_292;
assign r4_292 = in[3]? r3_584 : r3_583;
wire r4_293;
assign r4_293 = in[3]? r3_586 : r3_585;
wire r4_294;
assign r4_294 = in[3]? r3_588 : r3_587;
wire r4_295;
assign r4_295 = in[3]? r3_590 : r3_589;
wire r4_296;
assign r4_296 = in[3]? r3_592 : r3_591;
wire r4_297;
assign r4_297 = in[3]? r3_594 : r3_593;
wire r4_298;
assign r4_298 = in[3]? r3_596 : r3_595;
wire r4_299;
assign r4_299 = in[3]? r3_598 : r3_597;
wire r4_300;
assign r4_300 = in[3]? r3_600 : r3_599;
wire r4_301;
assign r4_301 = in[3]? r3_602 : r3_601;
wire r4_302;
assign r4_302 = in[3]? r3_604 : r3_603;
wire r4_303;
assign r4_303 = in[3]? r3_606 : r3_605;
wire r4_304;
assign r4_304 = in[3]? r3_608 : r3_607;
wire r4_305;
assign r4_305 = in[3]? r3_610 : r3_609;
wire r4_306;
assign r4_306 = in[3]? r3_612 : r3_611;
wire r4_307;
assign r4_307 = in[3]? r3_614 : r3_613;
wire r4_308;
assign r4_308 = in[3]? r3_616 : r3_615;
wire r4_309;
assign r4_309 = in[3]? r3_618 : r3_617;
wire r4_310;
assign r4_310 = in[3]? r3_620 : r3_619;
wire r4_311;
assign r4_311 = in[3]? r3_622 : r3_621;
wire r4_312;
assign r4_312 = in[3]? r3_624 : r3_623;
wire r4_313;
assign r4_313 = in[3]? r3_626 : r3_625;
wire r4_314;
assign r4_314 = in[3]? r3_628 : r3_627;
wire r4_315;
assign r4_315 = in[3]? r3_630 : r3_629;
wire r4_316;
assign r4_316 = in[3]? r3_632 : r3_631;
wire r4_317;
assign r4_317 = in[3]? r3_634 : r3_633;
wire r4_318;
assign r4_318 = in[3]? r3_636 : r3_635;
wire r4_319;
assign r4_319 = in[3]? r3_638 : r3_637;
wire r4_320;
assign r4_320 = in[3]? r3_640 : r3_639;
wire r4_321;
assign r4_321 = in[3]? r3_642 : r3_641;
wire r4_322;
assign r4_322 = in[3]? r3_644 : r3_643;
wire r4_323;
assign r4_323 = in[3]? r3_646 : r3_645;
wire r4_324;
assign r4_324 = in[3]? r3_648 : r3_647;
wire r4_325;
assign r4_325 = in[3]? r3_650 : r3_649;
wire r4_326;
assign r4_326 = in[3]? r3_652 : r3_651;
wire r4_327;
assign r4_327 = in[3]? r3_654 : r3_653;
wire r4_328;
assign r4_328 = in[3]? r3_656 : r3_655;
wire r4_329;
assign r4_329 = in[3]? r3_658 : r3_657;
wire r4_330;
assign r4_330 = in[3]? r3_660 : r3_659;
wire r4_331;
assign r4_331 = in[3]? r3_662 : r3_661;
wire r4_332;
assign r4_332 = in[3]? r3_664 : r3_663;
wire r4_333;
assign r4_333 = in[3]? r3_666 : r3_665;
wire r4_334;
assign r4_334 = in[3]? r3_668 : r3_667;
wire r4_335;
assign r4_335 = in[3]? r3_670 : r3_669;
wire r4_336;
assign r4_336 = in[3]? r3_672 : r3_671;
wire r4_337;
assign r4_337 = in[3]? r3_674 : r3_673;
wire r4_338;
assign r4_338 = in[3]? r3_676 : r3_675;
wire r4_339;
assign r4_339 = in[3]? r3_678 : r3_677;
wire r4_340;
assign r4_340 = in[3]? r3_680 : r3_679;
wire r4_341;
assign r4_341 = in[3]? r3_682 : r3_681;
wire r4_342;
assign r4_342 = in[3]? r3_684 : r3_683;
wire r4_343;
assign r4_343 = in[3]? r3_686 : r3_685;
wire r4_344;
assign r4_344 = in[3]? r3_688 : r3_687;
wire r4_345;
assign r4_345 = in[3]? r3_690 : r3_689;
wire r4_346;
assign r4_346 = in[3]? r3_692 : r3_691;
wire r4_347;
assign r4_347 = in[3]? r3_694 : r3_693;
wire r4_348;
assign r4_348 = in[3]? r3_696 : r3_695;
wire r4_349;
assign r4_349 = in[3]? r3_698 : r3_697;
wire r4_350;
assign r4_350 = in[3]? r3_700 : r3_699;
wire r4_351;
assign r4_351 = in[3]? r3_702 : r3_701;
wire r4_352;
assign r4_352 = in[3]? r3_704 : r3_703;
wire r4_353;
assign r4_353 = in[3]? r3_706 : r3_705;
wire r4_354;
assign r4_354 = in[3]? r3_708 : r3_707;
wire r4_355;
assign r4_355 = in[3]? r3_710 : r3_709;
wire r4_356;
assign r4_356 = in[3]? r3_712 : r3_711;
wire r4_357;
assign r4_357 = in[3]? r3_714 : r3_713;
wire r4_358;
assign r4_358 = in[3]? r3_716 : r3_715;
wire r4_359;
assign r4_359 = in[3]? r3_718 : r3_717;
wire r4_360;
assign r4_360 = in[3]? r3_720 : r3_719;
wire r4_361;
assign r4_361 = in[3]? r3_722 : r3_721;
wire r4_362;
assign r4_362 = in[3]? r3_724 : r3_723;
wire r4_363;
assign r4_363 = in[3]? r3_726 : r3_725;
wire r4_364;
assign r4_364 = in[3]? r3_728 : r3_727;
wire r4_365;
assign r4_365 = in[3]? r3_730 : r3_729;
wire r4_366;
assign r4_366 = in[3]? r3_732 : r3_731;
wire r4_367;
assign r4_367 = in[3]? r3_734 : r3_733;
wire r4_368;
assign r4_368 = in[3]? r3_736 : r3_735;
wire r4_369;
assign r4_369 = in[3]? r3_738 : r3_737;
wire r4_370;
assign r4_370 = in[3]? r3_740 : r3_739;
wire r4_371;
assign r4_371 = in[3]? r3_742 : r3_741;
wire r4_372;
assign r4_372 = in[3]? r3_744 : r3_743;
wire r4_373;
assign r4_373 = in[3]? r3_746 : r3_745;
wire r4_374;
assign r4_374 = in[3]? r3_748 : r3_747;
wire r4_375;
assign r4_375 = in[3]? r3_750 : r3_749;
wire r4_376;
assign r4_376 = in[3]? r3_752 : r3_751;
wire r4_377;
assign r4_377 = in[3]? r3_754 : r3_753;
wire r4_378;
assign r4_378 = in[3]? r3_756 : r3_755;
wire r4_379;
assign r4_379 = in[3]? r3_758 : r3_757;
wire r4_380;
assign r4_380 = in[3]? r3_760 : r3_759;
wire r4_381;
assign r4_381 = in[3]? r3_762 : r3_761;
wire r4_382;
assign r4_382 = in[3]? r3_764 : r3_763;
wire r4_383;
assign r4_383 = in[3]? r3_766 : r3_765;
wire r4_384;
assign r4_384 = in[3]? r3_768 : r3_767;
wire r4_385;
assign r4_385 = in[3]? r3_770 : r3_769;
wire r4_386;
assign r4_386 = in[3]? r3_772 : r3_771;
wire r4_387;
assign r4_387 = in[3]? r3_774 : r3_773;
wire r4_388;
assign r4_388 = in[3]? r3_776 : r3_775;
wire r4_389;
assign r4_389 = in[3]? r3_778 : r3_777;
wire r4_390;
assign r4_390 = in[3]? r3_780 : r3_779;
wire r4_391;
assign r4_391 = in[3]? r3_782 : r3_781;
wire r4_392;
assign r4_392 = in[3]? r3_784 : r3_783;
wire r4_393;
assign r4_393 = in[3]? r3_786 : r3_785;
wire r4_394;
assign r4_394 = in[3]? r3_788 : r3_787;
wire r4_395;
assign r4_395 = in[3]? r3_790 : r3_789;
wire r4_396;
assign r4_396 = in[3]? r3_792 : r3_791;
wire r4_397;
assign r4_397 = in[3]? r3_794 : r3_793;
wire r4_398;
assign r4_398 = in[3]? r3_796 : r3_795;
wire r4_399;
assign r4_399 = in[3]? r3_798 : r3_797;
wire r4_400;
assign r4_400 = in[3]? r3_800 : r3_799;
wire r4_401;
assign r4_401 = in[3]? r3_802 : r3_801;
wire r4_402;
assign r4_402 = in[3]? r3_804 : r3_803;
wire r4_403;
assign r4_403 = in[3]? r3_806 : r3_805;
wire r4_404;
assign r4_404 = in[3]? r3_808 : r3_807;
wire r4_405;
assign r4_405 = in[3]? r3_810 : r3_809;
wire r4_406;
assign r4_406 = in[3]? r3_812 : r3_811;
wire r4_407;
assign r4_407 = in[3]? r3_814 : r3_813;
wire r4_408;
assign r4_408 = in[3]? r3_816 : r3_815;
wire r4_409;
assign r4_409 = in[3]? r3_818 : r3_817;
wire r4_410;
assign r4_410 = in[3]? r3_820 : r3_819;
wire r4_411;
assign r4_411 = in[3]? r3_822 : r3_821;
wire r4_412;
assign r4_412 = in[3]? r3_824 : r3_823;
wire r4_413;
assign r4_413 = in[3]? r3_826 : r3_825;
wire r4_414;
assign r4_414 = in[3]? r3_828 : r3_827;
wire r4_415;
assign r4_415 = in[3]? r3_830 : r3_829;
wire r4_416;
assign r4_416 = in[3]? r3_832 : r3_831;
wire r4_417;
assign r4_417 = in[3]? r3_834 : r3_833;
wire r4_418;
assign r4_418 = in[3]? r3_836 : r3_835;
wire r4_419;
assign r4_419 = in[3]? r3_838 : r3_837;
wire r4_420;
assign r4_420 = in[3]? r3_840 : r3_839;
wire r4_421;
assign r4_421 = in[3]? r3_842 : r3_841;
wire r4_422;
assign r4_422 = in[3]? r3_844 : r3_843;
wire r4_423;
assign r4_423 = in[3]? r3_846 : r3_845;
wire r4_424;
assign r4_424 = in[3]? r3_848 : r3_847;
wire r4_425;
assign r4_425 = in[3]? r3_850 : r3_849;
wire r4_426;
assign r4_426 = in[3]? r3_852 : r3_851;
wire r4_427;
assign r4_427 = in[3]? r3_854 : r3_853;
wire r4_428;
assign r4_428 = in[3]? r3_856 : r3_855;
wire r4_429;
assign r4_429 = in[3]? r3_858 : r3_857;
wire r4_430;
assign r4_430 = in[3]? r3_860 : r3_859;
wire r4_431;
assign r4_431 = in[3]? r3_862 : r3_861;
wire r4_432;
assign r4_432 = in[3]? r3_864 : r3_863;
wire r4_433;
assign r4_433 = in[3]? r3_866 : r3_865;
wire r4_434;
assign r4_434 = in[3]? r3_868 : r3_867;
wire r4_435;
assign r4_435 = in[3]? r3_870 : r3_869;
wire r4_436;
assign r4_436 = in[3]? r3_872 : r3_871;
wire r4_437;
assign r4_437 = in[3]? r3_874 : r3_873;
wire r4_438;
assign r4_438 = in[3]? r3_876 : r3_875;
wire r4_439;
assign r4_439 = in[3]? r3_878 : r3_877;
wire r4_440;
assign r4_440 = in[3]? r3_880 : r3_879;
wire r4_441;
assign r4_441 = in[3]? r3_882 : r3_881;
wire r4_442;
assign r4_442 = in[3]? r3_884 : r3_883;
wire r4_443;
assign r4_443 = in[3]? r3_886 : r3_885;
wire r4_444;
assign r4_444 = in[3]? r3_888 : r3_887;
wire r4_445;
assign r4_445 = in[3]? r3_890 : r3_889;
wire r4_446;
assign r4_446 = in[3]? r3_892 : r3_891;
wire r4_447;
assign r4_447 = in[3]? r3_894 : r3_893;
wire r4_448;
assign r4_448 = in[3]? r3_896 : r3_895;
wire r4_449;
assign r4_449 = in[3]? r3_898 : r3_897;
wire r4_450;
assign r4_450 = in[3]? r3_900 : r3_899;
wire r4_451;
assign r4_451 = in[3]? r3_902 : r3_901;
wire r4_452;
assign r4_452 = in[3]? r3_904 : r3_903;
wire r4_453;
assign r4_453 = in[3]? r3_906 : r3_905;
wire r4_454;
assign r4_454 = in[3]? r3_908 : r3_907;
wire r4_455;
assign r4_455 = in[3]? r3_910 : r3_909;
wire r4_456;
assign r4_456 = in[3]? r3_912 : r3_911;
wire r4_457;
assign r4_457 = in[3]? r3_914 : r3_913;
wire r4_458;
assign r4_458 = in[3]? r3_916 : r3_915;
wire r4_459;
assign r4_459 = in[3]? r3_918 : r3_917;
wire r4_460;
assign r4_460 = in[3]? r3_920 : r3_919;
wire r4_461;
assign r4_461 = in[3]? r3_922 : r3_921;
wire r4_462;
assign r4_462 = in[3]? r3_924 : r3_923;
wire r4_463;
assign r4_463 = in[3]? r3_926 : r3_925;
wire r4_464;
assign r4_464 = in[3]? r3_928 : r3_927;
wire r4_465;
assign r4_465 = in[3]? r3_930 : r3_929;
wire r4_466;
assign r4_466 = in[3]? r3_932 : r3_931;
wire r4_467;
assign r4_467 = in[3]? r3_934 : r3_933;
wire r4_468;
assign r4_468 = in[3]? r3_936 : r3_935;
wire r4_469;
assign r4_469 = in[3]? r3_938 : r3_937;
wire r4_470;
assign r4_470 = in[3]? r3_940 : r3_939;
wire r4_471;
assign r4_471 = in[3]? r3_942 : r3_941;
wire r4_472;
assign r4_472 = in[3]? r3_944 : r3_943;
wire r4_473;
assign r4_473 = in[3]? r3_946 : r3_945;
wire r4_474;
assign r4_474 = in[3]? r3_948 : r3_947;
wire r4_475;
assign r4_475 = in[3]? r3_950 : r3_949;
wire r4_476;
assign r4_476 = in[3]? r3_952 : r3_951;
wire r4_477;
assign r4_477 = in[3]? r3_954 : r3_953;
wire r4_478;
assign r4_478 = in[3]? r3_956 : r3_955;
wire r4_479;
assign r4_479 = in[3]? r3_958 : r3_957;
wire r4_480;
assign r4_480 = in[3]? r3_960 : r3_959;
wire r4_481;
assign r4_481 = in[3]? r3_962 : r3_961;
wire r4_482;
assign r4_482 = in[3]? r3_964 : r3_963;
wire r4_483;
assign r4_483 = in[3]? r3_966 : r3_965;
wire r4_484;
assign r4_484 = in[3]? r3_968 : r3_967;
wire r4_485;
assign r4_485 = in[3]? r3_970 : r3_969;
wire r4_486;
assign r4_486 = in[3]? r3_972 : r3_971;
wire r4_487;
assign r4_487 = in[3]? r3_974 : r3_973;
wire r4_488;
assign r4_488 = in[3]? r3_976 : r3_975;
wire r4_489;
assign r4_489 = in[3]? r3_978 : r3_977;
wire r4_490;
assign r4_490 = in[3]? r3_980 : r3_979;
wire r4_491;
assign r4_491 = in[3]? r3_982 : r3_981;
wire r4_492;
assign r4_492 = in[3]? r3_984 : r3_983;
wire r4_493;
assign r4_493 = in[3]? r3_986 : r3_985;
wire r4_494;
assign r4_494 = in[3]? r3_988 : r3_987;
wire r4_495;
assign r4_495 = in[3]? r3_990 : r3_989;
wire r4_496;
assign r4_496 = in[3]? r3_992 : r3_991;
wire r4_497;
assign r4_497 = in[3]? r3_994 : r3_993;
wire r4_498;
assign r4_498 = in[3]? r3_996 : r3_995;
wire r4_499;
assign r4_499 = in[3]? r3_998 : r3_997;
wire r4_500;
assign r4_500 = in[3]? r3_1000 : r3_999;
wire r4_501;
assign r4_501 = in[3]? r3_1002 : r3_1001;
wire r4_502;
assign r4_502 = in[3]? r3_1004 : r3_1003;
wire r4_503;
assign r4_503 = in[3]? r3_1006 : r3_1005;
wire r4_504;
assign r4_504 = in[3]? r3_1008 : r3_1007;
wire r4_505;
assign r4_505 = in[3]? r3_1010 : r3_1009;
wire r4_506;
assign r4_506 = in[3]? r3_1012 : r3_1011;
wire r4_507;
assign r4_507 = in[3]? r3_1014 : r3_1013;
wire r4_508;
assign r4_508 = in[3]? r3_1016 : r3_1015;
wire r4_509;
assign r4_509 = in[3]? r3_1018 : r3_1017;
wire r4_510;
assign r4_510 = in[3]? r3_1020 : r3_1019;
wire r4_511;
assign r4_511 = in[3]? r3_1022 : r3_1021;
wire r4_512;
assign r4_512 = in[3]? r3_1024 : r3_1023;
wire r4_513;
assign r4_513 = in[3]? r3_1026 : r3_1025;
wire r4_514;
assign r4_514 = in[3]? r3_1028 : r3_1027;
wire r4_515;
assign r4_515 = in[3]? r3_1030 : r3_1029;
wire r4_516;
assign r4_516 = in[3]? r3_1032 : r3_1031;
wire r4_517;
assign r4_517 = in[3]? r3_1034 : r3_1033;
wire r4_518;
assign r4_518 = in[3]? r3_1036 : r3_1035;
wire r4_519;
assign r4_519 = in[3]? r3_1038 : r3_1037;
wire r4_520;
assign r4_520 = in[3]? r3_1040 : r3_1039;
wire r4_521;
assign r4_521 = in[3]? r3_1042 : r3_1041;
wire r4_522;
assign r4_522 = in[3]? r3_1044 : r3_1043;
wire r4_523;
assign r4_523 = in[3]? r3_1046 : r3_1045;
wire r4_524;
assign r4_524 = in[3]? r3_1048 : r3_1047;
wire r4_525;
assign r4_525 = in[3]? r3_1050 : r3_1049;
wire r4_526;
assign r4_526 = in[3]? r3_1052 : r3_1051;
wire r4_527;
assign r4_527 = in[3]? r3_1054 : r3_1053;
wire r4_528;
assign r4_528 = in[3]? r3_1056 : r3_1055;
wire r4_529;
assign r4_529 = in[3]? r3_1058 : r3_1057;
wire r4_530;
assign r4_530 = in[3]? r3_1060 : r3_1059;
wire r4_531;
assign r4_531 = in[3]? r3_1062 : r3_1061;
wire r4_532;
assign r4_532 = in[3]? r3_1064 : r3_1063;
wire r4_533;
assign r4_533 = in[3]? r3_1066 : r3_1065;
wire r4_534;
assign r4_534 = in[3]? r3_1068 : r3_1067;
wire r4_535;
assign r4_535 = in[3]? r3_1070 : r3_1069;
wire r4_536;
assign r4_536 = in[3]? r3_1072 : r3_1071;
wire r4_537;
assign r4_537 = in[3]? r3_1074 : r3_1073;
wire r4_538;
assign r4_538 = in[3]? r3_1076 : r3_1075;
wire r4_539;
assign r4_539 = in[3]? r3_1078 : r3_1077;
wire r4_540;
assign r4_540 = in[3]? r3_1080 : r3_1079;
wire r4_541;
assign r4_541 = in[3]? r3_1082 : r3_1081;
wire r4_542;
assign r4_542 = in[3]? r3_1084 : r3_1083;
wire r4_543;
assign r4_543 = in[3]? r3_1086 : r3_1085;
wire r4_544;
assign r4_544 = in[3]? r3_1088 : r3_1087;
wire r4_545;
assign r4_545 = in[3]? r3_1090 : r3_1089;
wire r4_546;
assign r4_546 = in[3]? r3_1092 : r3_1091;
wire r4_547;
assign r4_547 = in[3]? r3_1094 : r3_1093;
wire r4_548;
assign r4_548 = in[3]? r3_1096 : r3_1095;
wire r4_549;
assign r4_549 = in[3]? r3_1098 : r3_1097;
wire r4_550;
assign r4_550 = in[3]? r3_1100 : r3_1099;
wire r4_551;
assign r4_551 = in[3]? r3_1102 : r3_1101;
wire r4_552;
assign r4_552 = in[3]? r3_1104 : r3_1103;
wire r4_553;
assign r4_553 = in[3]? r3_1106 : r3_1105;
wire r4_554;
assign r4_554 = in[3]? r3_1108 : r3_1107;
wire r4_555;
assign r4_555 = in[3]? r3_1110 : r3_1109;
wire r4_556;
assign r4_556 = in[3]? r3_1112 : r3_1111;
wire r4_557;
assign r4_557 = in[3]? r3_1114 : r3_1113;
wire r4_558;
assign r4_558 = in[3]? r3_1116 : r3_1115;
wire r4_559;
assign r4_559 = in[3]? r3_1118 : r3_1117;
wire r4_560;
assign r4_560 = in[3]? r3_1120 : r3_1119;
wire r4_561;
assign r4_561 = in[3]? r3_1122 : r3_1121;
wire r4_562;
assign r4_562 = in[3]? r3_1124 : r3_1123;
wire r4_563;
assign r4_563 = in[3]? r3_1126 : r3_1125;
wire r4_564;
assign r4_564 = in[3]? r3_1128 : r3_1127;
wire r4_565;
assign r4_565 = in[3]? r3_1130 : r3_1129;
wire r4_566;
assign r4_566 = in[3]? r3_1132 : r3_1131;
wire r4_567;
assign r4_567 = in[3]? r3_1134 : r3_1133;
wire r4_568;
assign r4_568 = in[3]? r3_1136 : r3_1135;
wire r4_569;
assign r4_569 = in[3]? r3_1138 : r3_1137;
wire r4_570;
assign r4_570 = in[3]? r3_1140 : r3_1139;
wire r4_571;
assign r4_571 = in[3]? r3_1142 : r3_1141;
wire r4_572;
assign r4_572 = in[3]? r3_1144 : r3_1143;
wire r4_573;
assign r4_573 = in[3]? r3_1146 : r3_1145;
wire r4_574;
assign r4_574 = in[3]? r3_1148 : r3_1147;
wire r4_575;
assign r4_575 = in[3]? r3_1150 : r3_1149;
wire r4_576;
assign r4_576 = in[3]? r3_1152 : r3_1151;
wire r4_577;
assign r4_577 = in[3]? r3_1154 : r3_1153;
wire r4_578;
assign r4_578 = in[3]? r3_1156 : r3_1155;
wire r4_579;
assign r4_579 = in[3]? r3_1158 : r3_1157;
wire r4_580;
assign r4_580 = in[3]? r3_1160 : r3_1159;
wire r4_581;
assign r4_581 = in[3]? r3_1162 : r3_1161;
wire r4_582;
assign r4_582 = in[3]? r3_1164 : r3_1163;
wire r4_583;
assign r4_583 = in[3]? r3_1166 : r3_1165;
wire r4_584;
assign r4_584 = in[3]? r3_1168 : r3_1167;
wire r4_585;
assign r4_585 = in[3]? r3_1170 : r3_1169;
wire r4_586;
assign r4_586 = in[3]? r3_1172 : r3_1171;
wire r4_587;
assign r4_587 = in[3]? r3_1174 : r3_1173;
wire r4_588;
assign r4_588 = in[3]? r3_1176 : r3_1175;
wire r4_589;
assign r4_589 = in[3]? r3_1178 : r3_1177;
wire r4_590;
assign r4_590 = in[3]? r3_1180 : r3_1179;
wire r4_591;
assign r4_591 = in[3]? r3_1182 : r3_1181;
wire r4_592;
assign r4_592 = in[3]? r3_1184 : r3_1183;
wire r4_593;
assign r4_593 = in[3]? r3_1186 : r3_1185;
wire r4_594;
assign r4_594 = in[3]? r3_1188 : r3_1187;
wire r4_595;
assign r4_595 = in[3]? r3_1190 : r3_1189;
wire r4_596;
assign r4_596 = in[3]? r3_1192 : r3_1191;
wire r4_597;
assign r4_597 = in[3]? r3_1194 : r3_1193;
wire r4_598;
assign r4_598 = in[3]? r3_1196 : r3_1195;
wire r4_599;
assign r4_599 = in[3]? r3_1198 : r3_1197;
wire r4_600;
assign r4_600 = in[3]? r3_1200 : r3_1199;
wire r4_601;
assign r4_601 = in[3]? r3_1202 : r3_1201;
wire r4_602;
assign r4_602 = in[3]? r3_1204 : r3_1203;
wire r4_603;
assign r4_603 = in[3]? r3_1206 : r3_1205;
wire r4_604;
assign r4_604 = in[3]? r3_1208 : r3_1207;
wire r4_605;
assign r4_605 = in[3]? r3_1210 : r3_1209;
wire r4_606;
assign r4_606 = in[3]? r3_1212 : r3_1211;
wire r4_607;
assign r4_607 = in[3]? r3_1214 : r3_1213;
wire r4_608;
assign r4_608 = in[3]? r3_1216 : r3_1215;
wire r4_609;
assign r4_609 = in[3]? r3_1218 : r3_1217;
wire r4_610;
assign r4_610 = in[3]? r3_1220 : r3_1219;
wire r4_611;
assign r4_611 = in[3]? r3_1222 : r3_1221;
wire r4_612;
assign r4_612 = in[3]? r3_1224 : r3_1223;
wire r4_613;
assign r4_613 = in[3]? r3_1226 : r3_1225;
wire r4_614;
assign r4_614 = in[3]? r3_1228 : r3_1227;
wire r4_615;
assign r4_615 = in[3]? r3_1230 : r3_1229;
wire r4_616;
assign r4_616 = in[3]? r3_1232 : r3_1231;
wire r4_617;
assign r4_617 = in[3]? r3_1234 : r3_1233;
wire r4_618;
assign r4_618 = in[3]? r3_1236 : r3_1235;
wire r4_619;
assign r4_619 = in[3]? r3_1238 : r3_1237;
wire r4_620;
assign r4_620 = in[3]? r3_1240 : r3_1239;
wire r4_621;
assign r4_621 = in[3]? r3_1242 : r3_1241;
wire r4_622;
assign r4_622 = in[3]? r3_1244 : r3_1243;
wire r4_623;
assign r4_623 = in[3]? r3_1246 : r3_1245;
wire r4_624;
assign r4_624 = in[3]? r3_1248 : r3_1247;
wire r4_625;
assign r4_625 = in[3]? r3_1250 : r3_1249;
wire r4_626;
assign r4_626 = in[3]? r3_1252 : r3_1251;
wire r4_627;
assign r4_627 = in[3]? r3_1254 : r3_1253;
wire r4_628;
assign r4_628 = in[3]? r3_1256 : r3_1255;
wire r4_629;
assign r4_629 = in[3]? r3_1258 : r3_1257;
wire r4_630;
assign r4_630 = in[3]? r3_1260 : r3_1259;
wire r4_631;
assign r4_631 = in[3]? r3_1262 : r3_1261;
wire r4_632;
assign r4_632 = in[3]? r3_1264 : r3_1263;
wire r4_633;
assign r4_633 = in[3]? r3_1266 : r3_1265;
wire r4_634;
assign r4_634 = in[3]? r3_1268 : r3_1267;
wire r4_635;
assign r4_635 = in[3]? r3_1270 : r3_1269;
wire r4_636;
assign r4_636 = in[3]? r3_1272 : r3_1271;
wire r4_637;
assign r4_637 = in[3]? r3_1274 : r3_1273;
wire r4_638;
assign r4_638 = in[3]? r3_1276 : r3_1275;
wire r4_639;
assign r4_639 = in[3]? r3_1278 : r3_1277;
wire r4_640;
assign r4_640 = in[3]? r3_1280 : r3_1279;
wire r4_641;
assign r4_641 = in[3]? r3_1282 : r3_1281;
wire r4_642;
assign r4_642 = in[3]? r3_1284 : r3_1283;
wire r4_643;
assign r4_643 = in[3]? r3_1286 : r3_1285;
wire r4_644;
assign r4_644 = in[3]? r3_1288 : r3_1287;
wire r4_645;
assign r4_645 = in[3]? r3_1290 : r3_1289;
wire r4_646;
assign r4_646 = in[3]? r3_1292 : r3_1291;
wire r4_647;
assign r4_647 = in[3]? r3_1294 : r3_1293;
wire r4_648;
assign r4_648 = in[3]? r3_1296 : r3_1295;
wire r4_649;
assign r4_649 = in[3]? r3_1298 : r3_1297;
wire r4_650;
assign r4_650 = in[3]? r3_1300 : r3_1299;
wire r4_651;
assign r4_651 = in[3]? r3_1302 : r3_1301;
wire r4_652;
assign r4_652 = in[3]? r3_1304 : r3_1303;
wire r4_653;
assign r4_653 = in[3]? r3_1306 : r3_1305;
wire r4_654;
assign r4_654 = in[3]? r3_1308 : r3_1307;
wire r4_655;
assign r4_655 = in[3]? r3_1310 : r3_1309;
wire r4_656;
assign r4_656 = in[3]? r3_1312 : r3_1311;
wire r4_657;
assign r4_657 = in[3]? r3_1314 : r3_1313;
wire r4_658;
assign r4_658 = in[3]? r3_1316 : r3_1315;
wire r4_659;
assign r4_659 = in[3]? r3_1318 : r3_1317;
wire r4_660;
assign r4_660 = in[3]? r3_1320 : r3_1319;
wire r4_661;
assign r4_661 = in[3]? r3_1322 : r3_1321;
wire r4_662;
assign r4_662 = in[3]? r3_1324 : r3_1323;
wire r4_663;
assign r4_663 = in[3]? r3_1326 : r3_1325;
wire r4_664;
assign r4_664 = in[3]? r3_1328 : r3_1327;
wire r4_665;
assign r4_665 = in[3]? r3_1330 : r3_1329;
wire r4_666;
assign r4_666 = in[3]? r3_1332 : r3_1331;
wire r4_667;
assign r4_667 = in[3]? r3_1334 : r3_1333;
wire r4_668;
assign r4_668 = in[3]? r3_1336 : r3_1335;
wire r4_669;
assign r4_669 = in[3]? r3_1338 : r3_1337;
wire r4_670;
assign r4_670 = in[3]? r3_1340 : r3_1339;
wire r4_671;
assign r4_671 = in[3]? r3_1342 : r3_1341;
wire r4_672;
assign r4_672 = in[3]? r3_1344 : r3_1343;
wire r4_673;
assign r4_673 = in[3]? r3_1346 : r3_1345;
wire r4_674;
assign r4_674 = in[3]? r3_1348 : r3_1347;
wire r4_675;
assign r4_675 = in[3]? r3_1350 : r3_1349;
wire r4_676;
assign r4_676 = in[3]? r3_1352 : r3_1351;
wire r4_677;
assign r4_677 = in[3]? r3_1354 : r3_1353;
wire r4_678;
assign r4_678 = in[3]? r3_1356 : r3_1355;
wire r4_679;
assign r4_679 = in[3]? r3_1358 : r3_1357;
wire r4_680;
assign r4_680 = in[3]? r3_1360 : r3_1359;
wire r4_681;
assign r4_681 = in[3]? r3_1362 : r3_1361;
wire r4_682;
assign r4_682 = in[3]? r3_1364 : r3_1363;
wire r4_683;
assign r4_683 = in[3]? r3_1366 : r3_1365;
wire r4_684;
assign r4_684 = in[3]? r3_1368 : r3_1367;
wire r4_685;
assign r4_685 = in[3]? r3_1370 : r3_1369;
wire r4_686;
assign r4_686 = in[3]? r3_1372 : r3_1371;
wire r4_687;
assign r4_687 = in[3]? r3_1374 : r3_1373;
wire r4_688;
assign r4_688 = in[3]? r3_1376 : r3_1375;
wire r4_689;
assign r4_689 = in[3]? r3_1378 : r3_1377;
wire r4_690;
assign r4_690 = in[3]? r3_1380 : r3_1379;
wire r4_691;
assign r4_691 = in[3]? r3_1382 : r3_1381;
wire r4_692;
assign r4_692 = in[3]? r3_1384 : r3_1383;
wire r4_693;
assign r4_693 = in[3]? r3_1386 : r3_1385;
wire r4_694;
assign r4_694 = in[3]? r3_1388 : r3_1387;
wire r4_695;
assign r4_695 = in[3]? r3_1390 : r3_1389;
wire r4_696;
assign r4_696 = in[3]? r3_1392 : r3_1391;
wire r4_697;
assign r4_697 = in[3]? r3_1394 : r3_1393;
wire r4_698;
assign r4_698 = in[3]? r3_1396 : r3_1395;
wire r4_699;
assign r4_699 = in[3]? r3_1398 : r3_1397;
wire r4_700;
assign r4_700 = in[3]? r3_1400 : r3_1399;
wire r4_701;
assign r4_701 = in[3]? r3_1402 : r3_1401;
wire r4_702;
assign r4_702 = in[3]? r3_1404 : r3_1403;
wire r4_703;
assign r4_703 = in[3]? r3_1406 : r3_1405;
wire r4_704;
assign r4_704 = in[3]? r3_1408 : r3_1407;
wire r4_705;
assign r4_705 = in[3]? r3_1410 : r3_1409;
wire r4_706;
assign r4_706 = in[3]? r3_1412 : r3_1411;
wire r4_707;
assign r4_707 = in[3]? r3_1414 : r3_1413;
wire r4_708;
assign r4_708 = in[3]? r3_1416 : r3_1415;
wire r4_709;
assign r4_709 = in[3]? r3_1418 : r3_1417;
wire r4_710;
assign r4_710 = in[3]? r3_1420 : r3_1419;
wire r4_711;
assign r4_711 = in[3]? r3_1422 : r3_1421;
wire r4_712;
assign r4_712 = in[3]? r3_1424 : r3_1423;
wire r4_713;
assign r4_713 = in[3]? r3_1426 : r3_1425;
wire r4_714;
assign r4_714 = in[3]? r3_1428 : r3_1427;
wire r4_715;
assign r4_715 = in[3]? r3_1430 : r3_1429;
wire r4_716;
assign r4_716 = in[3]? r3_1432 : r3_1431;
wire r4_717;
assign r4_717 = in[3]? r3_1434 : r3_1433;
wire r4_718;
assign r4_718 = in[3]? r3_1436 : r3_1435;
wire r4_719;
assign r4_719 = in[3]? r3_1438 : r3_1437;
wire r4_720;
assign r4_720 = in[3]? r3_1440 : r3_1439;
wire r4_721;
assign r4_721 = in[3]? r3_1442 : r3_1441;
wire r4_722;
assign r4_722 = in[3]? r3_1444 : r3_1443;
wire r4_723;
assign r4_723 = in[3]? r3_1446 : r3_1445;
wire r4_724;
assign r4_724 = in[3]? r3_1448 : r3_1447;
wire r4_725;
assign r4_725 = in[3]? r3_1450 : r3_1449;
wire r4_726;
assign r4_726 = in[3]? r3_1452 : r3_1451;
wire r4_727;
assign r4_727 = in[3]? r3_1454 : r3_1453;
wire r4_728;
assign r4_728 = in[3]? r3_1456 : r3_1455;
wire r4_729;
assign r4_729 = in[3]? r3_1458 : r3_1457;
wire r4_730;
assign r4_730 = in[3]? r3_1460 : r3_1459;
wire r4_731;
assign r4_731 = in[3]? r3_1462 : r3_1461;
wire r4_732;
assign r4_732 = in[3]? r3_1464 : r3_1463;
wire r4_733;
assign r4_733 = in[3]? r3_1466 : r3_1465;
wire r4_734;
assign r4_734 = in[3]? r3_1468 : r3_1467;
wire r4_735;
assign r4_735 = in[3]? r3_1470 : r3_1469;
wire r4_736;
assign r4_736 = in[3]? r3_1472 : r3_1471;
wire r4_737;
assign r4_737 = in[3]? r3_1474 : r3_1473;
wire r4_738;
assign r4_738 = in[3]? r3_1476 : r3_1475;
wire r4_739;
assign r4_739 = in[3]? r3_1478 : r3_1477;
wire r4_740;
assign r4_740 = in[3]? r3_1480 : r3_1479;
wire r4_741;
assign r4_741 = in[3]? r3_1482 : r3_1481;
wire r4_742;
assign r4_742 = in[3]? r3_1484 : r3_1483;
wire r4_743;
assign r4_743 = in[3]? r3_1486 : r3_1485;
wire r4_744;
assign r4_744 = in[3]? r3_1488 : r3_1487;
wire r4_745;
assign r4_745 = in[3]? r3_1490 : r3_1489;
wire r4_746;
assign r4_746 = in[3]? r3_1492 : r3_1491;
wire r4_747;
assign r4_747 = in[3]? r3_1494 : r3_1493;
wire r4_748;
assign r4_748 = in[3]? r3_1496 : r3_1495;
wire r4_749;
assign r4_749 = in[3]? r3_1498 : r3_1497;
wire r4_750;
assign r4_750 = in[3]? r3_1500 : r3_1499;
wire r4_751;
assign r4_751 = in[3]? r3_1502 : r3_1501;
wire r4_752;
assign r4_752 = in[3]? r3_1504 : r3_1503;
wire r4_753;
assign r4_753 = in[3]? r3_1506 : r3_1505;
wire r4_754;
assign r4_754 = in[3]? r3_1508 : r3_1507;
wire r4_755;
assign r4_755 = in[3]? r3_1510 : r3_1509;
wire r4_756;
assign r4_756 = in[3]? r3_1512 : r3_1511;
wire r4_757;
assign r4_757 = in[3]? r3_1514 : r3_1513;
wire r4_758;
assign r4_758 = in[3]? r3_1516 : r3_1515;
wire r4_759;
assign r4_759 = in[3]? r3_1518 : r3_1517;
wire r4_760;
assign r4_760 = in[3]? r3_1520 : r3_1519;
wire r4_761;
assign r4_761 = in[3]? r3_1522 : r3_1521;
wire r4_762;
assign r4_762 = in[3]? r3_1524 : r3_1523;
wire r4_763;
assign r4_763 = in[3]? r3_1526 : r3_1525;
wire r4_764;
assign r4_764 = in[3]? r3_1528 : r3_1527;
wire r4_765;
assign r4_765 = in[3]? r3_1530 : r3_1529;
wire r4_766;
assign r4_766 = in[3]? r3_1532 : r3_1531;
wire r4_767;
assign r4_767 = in[3]? r3_1534 : r3_1533;
wire r4_768;
assign r4_768 = in[3]? r3_1536 : r3_1535;
wire r4_769;
assign r4_769 = in[3]? r3_1538 : r3_1537;
wire r4_770;
assign r4_770 = in[3]? r3_1540 : r3_1539;
wire r4_771;
assign r4_771 = in[3]? r3_1542 : r3_1541;
wire r4_772;
assign r4_772 = in[3]? r3_1544 : r3_1543;
wire r4_773;
assign r4_773 = in[3]? r3_1546 : r3_1545;
wire r4_774;
assign r4_774 = in[3]? r3_1548 : r3_1547;
wire r4_775;
assign r4_775 = in[3]? r3_1550 : r3_1549;
wire r4_776;
assign r4_776 = in[3]? r3_1552 : r3_1551;
wire r4_777;
assign r4_777 = in[3]? r3_1554 : r3_1553;
wire r4_778;
assign r4_778 = in[3]? r3_1556 : r3_1555;
wire r4_779;
assign r4_779 = in[3]? r3_1558 : r3_1557;
wire r4_780;
assign r4_780 = in[3]? r3_1560 : r3_1559;
wire r4_781;
assign r4_781 = in[3]? r3_1562 : r3_1561;
wire r4_782;
assign r4_782 = in[3]? r3_1564 : r3_1563;
wire r4_783;
assign r4_783 = in[3]? r3_1566 : r3_1565;
wire r4_784;
assign r4_784 = in[3]? r3_1568 : r3_1567;
wire r4_785;
assign r4_785 = in[3]? r3_1570 : r3_1569;
wire r4_786;
assign r4_786 = in[3]? r3_1572 : r3_1571;
wire r4_787;
assign r4_787 = in[3]? r3_1574 : r3_1573;
wire r4_788;
assign r4_788 = in[3]? r3_1576 : r3_1575;
wire r4_789;
assign r4_789 = in[3]? r3_1578 : r3_1577;
wire r4_790;
assign r4_790 = in[3]? r3_1580 : r3_1579;
wire r4_791;
assign r4_791 = in[3]? r3_1582 : r3_1581;
wire r4_792;
assign r4_792 = in[3]? r3_1584 : r3_1583;
wire r4_793;
assign r4_793 = in[3]? r3_1586 : r3_1585;
wire r4_794;
assign r4_794 = in[3]? r3_1588 : r3_1587;
wire r4_795;
assign r4_795 = in[3]? r3_1590 : r3_1589;
wire r4_796;
assign r4_796 = in[3]? r3_1592 : r3_1591;
wire r4_797;
assign r4_797 = in[3]? r3_1594 : r3_1593;
wire r4_798;
assign r4_798 = in[3]? r3_1596 : r3_1595;
wire r4_799;
assign r4_799 = in[3]? r3_1598 : r3_1597;
wire r4_800;
assign r4_800 = in[3]? r3_1600 : r3_1599;
wire r4_801;
assign r4_801 = in[3]? r3_1602 : r3_1601;
wire r4_802;
assign r4_802 = in[3]? r3_1604 : r3_1603;
wire r4_803;
assign r4_803 = in[3]? r3_1606 : r3_1605;
wire r4_804;
assign r4_804 = in[3]? r3_1608 : r3_1607;
wire r4_805;
assign r4_805 = in[3]? r3_1610 : r3_1609;
wire r4_806;
assign r4_806 = in[3]? r3_1612 : r3_1611;
wire r4_807;
assign r4_807 = in[3]? r3_1614 : r3_1613;
wire r4_808;
assign r4_808 = in[3]? r3_1616 : r3_1615;
wire r4_809;
assign r4_809 = in[3]? r3_1618 : r3_1617;
wire r4_810;
assign r4_810 = in[3]? r3_1620 : r3_1619;
wire r4_811;
assign r4_811 = in[3]? r3_1622 : r3_1621;
wire r4_812;
assign r4_812 = in[3]? r3_1624 : r3_1623;
wire r4_813;
assign r4_813 = in[3]? r3_1626 : r3_1625;
wire r4_814;
assign r4_814 = in[3]? r3_1628 : r3_1627;
wire r4_815;
assign r4_815 = in[3]? r3_1630 : r3_1629;
wire r4_816;
assign r4_816 = in[3]? r3_1632 : r3_1631;
wire r4_817;
assign r4_817 = in[3]? r3_1634 : r3_1633;
wire r4_818;
assign r4_818 = in[3]? r3_1636 : r3_1635;
wire r4_819;
assign r4_819 = in[3]? r3_1638 : r3_1637;
wire r4_820;
assign r4_820 = in[3]? r3_1640 : r3_1639;
wire r4_821;
assign r4_821 = in[3]? r3_1642 : r3_1641;
wire r4_822;
assign r4_822 = in[3]? r3_1644 : r3_1643;
wire r4_823;
assign r4_823 = in[3]? r3_1646 : r3_1645;
wire r4_824;
assign r4_824 = in[3]? r3_1648 : r3_1647;
wire r4_825;
assign r4_825 = in[3]? r3_1650 : r3_1649;
wire r4_826;
assign r4_826 = in[3]? r3_1652 : r3_1651;
wire r4_827;
assign r4_827 = in[3]? r3_1654 : r3_1653;
wire r4_828;
assign r4_828 = in[3]? r3_1656 : r3_1655;
wire r4_829;
assign r4_829 = in[3]? r3_1658 : r3_1657;
wire r4_830;
assign r4_830 = in[3]? r3_1660 : r3_1659;
wire r4_831;
assign r4_831 = in[3]? r3_1662 : r3_1661;
wire r4_832;
assign r4_832 = in[3]? r3_1664 : r3_1663;
wire r4_833;
assign r4_833 = in[3]? r3_1666 : r3_1665;
wire r4_834;
assign r4_834 = in[3]? r3_1668 : r3_1667;
wire r4_835;
assign r4_835 = in[3]? r3_1670 : r3_1669;
wire r4_836;
assign r4_836 = in[3]? r3_1672 : r3_1671;
wire r4_837;
assign r4_837 = in[3]? r3_1674 : r3_1673;
wire r4_838;
assign r4_838 = in[3]? r3_1676 : r3_1675;
wire r4_839;
assign r4_839 = in[3]? r3_1678 : r3_1677;
wire r4_840;
assign r4_840 = in[3]? r3_1680 : r3_1679;
wire r4_841;
assign r4_841 = in[3]? r3_1682 : r3_1681;
wire r4_842;
assign r4_842 = in[3]? r3_1684 : r3_1683;
wire r4_843;
assign r4_843 = in[3]? r3_1686 : r3_1685;
wire r4_844;
assign r4_844 = in[3]? r3_1688 : r3_1687;
wire r4_845;
assign r4_845 = in[3]? r3_1690 : r3_1689;
wire r4_846;
assign r4_846 = in[3]? r3_1692 : r3_1691;
wire r4_847;
assign r4_847 = in[3]? r3_1694 : r3_1693;
wire r4_848;
assign r4_848 = in[3]? r3_1696 : r3_1695;
wire r4_849;
assign r4_849 = in[3]? r3_1698 : r3_1697;
wire r4_850;
assign r4_850 = in[3]? r3_1700 : r3_1699;
wire r4_851;
assign r4_851 = in[3]? r3_1702 : r3_1701;
wire r4_852;
assign r4_852 = in[3]? r3_1704 : r3_1703;
wire r4_853;
assign r4_853 = in[3]? r3_1706 : r3_1705;
wire r4_854;
assign r4_854 = in[3]? r3_1708 : r3_1707;
wire r4_855;
assign r4_855 = in[3]? r3_1710 : r3_1709;
wire r4_856;
assign r4_856 = in[3]? r3_1712 : r3_1711;
wire r4_857;
assign r4_857 = in[3]? r3_1714 : r3_1713;
wire r4_858;
assign r4_858 = in[3]? r3_1716 : r3_1715;
wire r4_859;
assign r4_859 = in[3]? r3_1718 : r3_1717;
wire r4_860;
assign r4_860 = in[3]? r3_1720 : r3_1719;
wire r4_861;
assign r4_861 = in[3]? r3_1722 : r3_1721;
wire r4_862;
assign r4_862 = in[3]? r3_1724 : r3_1723;
wire r4_863;
assign r4_863 = in[3]? r3_1726 : r3_1725;
wire r4_864;
assign r4_864 = in[3]? r3_1728 : r3_1727;
wire r4_865;
assign r4_865 = in[3]? r3_1730 : r3_1729;
wire r4_866;
assign r4_866 = in[3]? r3_1732 : r3_1731;
wire r4_867;
assign r4_867 = in[3]? r3_1734 : r3_1733;
wire r4_868;
assign r4_868 = in[3]? r3_1736 : r3_1735;
wire r4_869;
assign r4_869 = in[3]? r3_1738 : r3_1737;
wire r4_870;
assign r4_870 = in[3]? r3_1740 : r3_1739;
wire r4_871;
assign r4_871 = in[3]? r3_1742 : r3_1741;
wire r4_872;
assign r4_872 = in[3]? r3_1744 : r3_1743;
wire r4_873;
assign r4_873 = in[3]? r3_1746 : r3_1745;
wire r4_874;
assign r4_874 = in[3]? r3_1748 : r3_1747;
wire r4_875;
assign r4_875 = in[3]? r3_1750 : r3_1749;
wire r4_876;
assign r4_876 = in[3]? r3_1752 : r3_1751;
wire r4_877;
assign r4_877 = in[3]? r3_1754 : r3_1753;
wire r4_878;
assign r4_878 = in[3]? r3_1756 : r3_1755;
wire r4_879;
assign r4_879 = in[3]? r3_1758 : r3_1757;
wire r4_880;
assign r4_880 = in[3]? r3_1760 : r3_1759;
wire r4_881;
assign r4_881 = in[3]? r3_1762 : r3_1761;
wire r4_882;
assign r4_882 = in[3]? r3_1764 : r3_1763;
wire r4_883;
assign r4_883 = in[3]? r3_1766 : r3_1765;
wire r4_884;
assign r4_884 = in[3]? r3_1768 : r3_1767;
wire r4_885;
assign r4_885 = in[3]? r3_1770 : r3_1769;
wire r4_886;
assign r4_886 = in[3]? r3_1772 : r3_1771;
wire r4_887;
assign r4_887 = in[3]? r3_1774 : r3_1773;
wire r4_888;
assign r4_888 = in[3]? r3_1776 : r3_1775;
wire r4_889;
assign r4_889 = in[3]? r3_1778 : r3_1777;
wire r4_890;
assign r4_890 = in[3]? r3_1780 : r3_1779;
wire r4_891;
assign r4_891 = in[3]? r3_1782 : r3_1781;
wire r4_892;
assign r4_892 = in[3]? r3_1784 : r3_1783;
wire r4_893;
assign r4_893 = in[3]? r3_1786 : r3_1785;
wire r4_894;
assign r4_894 = in[3]? r3_1788 : r3_1787;
wire r4_895;
assign r4_895 = in[3]? r3_1790 : r3_1789;
wire r4_896;
assign r4_896 = in[3]? r3_1792 : r3_1791;
wire r4_897;
assign r4_897 = in[3]? r3_1794 : r3_1793;
wire r4_898;
assign r4_898 = in[3]? r3_1796 : r3_1795;
wire r4_899;
assign r4_899 = in[3]? r3_1798 : r3_1797;
wire r4_900;
assign r4_900 = in[3]? r3_1800 : r3_1799;
wire r4_901;
assign r4_901 = in[3]? r3_1802 : r3_1801;
wire r4_902;
assign r4_902 = in[3]? r3_1804 : r3_1803;
wire r4_903;
assign r4_903 = in[3]? r3_1806 : r3_1805;
wire r4_904;
assign r4_904 = in[3]? r3_1808 : r3_1807;
wire r4_905;
assign r4_905 = in[3]? r3_1810 : r3_1809;
wire r4_906;
assign r4_906 = in[3]? r3_1812 : r3_1811;
wire r4_907;
assign r4_907 = in[3]? r3_1814 : r3_1813;
wire r4_908;
assign r4_908 = in[3]? r3_1816 : r3_1815;
wire r4_909;
assign r4_909 = in[3]? r3_1818 : r3_1817;
wire r4_910;
assign r4_910 = in[3]? r3_1820 : r3_1819;
wire r4_911;
assign r4_911 = in[3]? r3_1822 : r3_1821;
wire r4_912;
assign r4_912 = in[3]? r3_1824 : r3_1823;
wire r4_913;
assign r4_913 = in[3]? r3_1826 : r3_1825;
wire r4_914;
assign r4_914 = in[3]? r3_1828 : r3_1827;
wire r4_915;
assign r4_915 = in[3]? r3_1830 : r3_1829;
wire r4_916;
assign r4_916 = in[3]? r3_1832 : r3_1831;
wire r4_917;
assign r4_917 = in[3]? r3_1834 : r3_1833;
wire r4_918;
assign r4_918 = in[3]? r3_1836 : r3_1835;
wire r4_919;
assign r4_919 = in[3]? r3_1838 : r3_1837;
wire r4_920;
assign r4_920 = in[3]? r3_1840 : r3_1839;
wire r4_921;
assign r4_921 = in[3]? r3_1842 : r3_1841;
wire r4_922;
assign r4_922 = in[3]? r3_1844 : r3_1843;
wire r4_923;
assign r4_923 = in[3]? r3_1846 : r3_1845;
wire r4_924;
assign r4_924 = in[3]? r3_1848 : r3_1847;
wire r4_925;
assign r4_925 = in[3]? r3_1850 : r3_1849;
wire r4_926;
assign r4_926 = in[3]? r3_1852 : r3_1851;
wire r4_927;
assign r4_927 = in[3]? r3_1854 : r3_1853;
wire r4_928;
assign r4_928 = in[3]? r3_1856 : r3_1855;
wire r4_929;
assign r4_929 = in[3]? r3_1858 : r3_1857;
wire r4_930;
assign r4_930 = in[3]? r3_1860 : r3_1859;
wire r4_931;
assign r4_931 = in[3]? r3_1862 : r3_1861;
wire r4_932;
assign r4_932 = in[3]? r3_1864 : r3_1863;
wire r4_933;
assign r4_933 = in[3]? r3_1866 : r3_1865;
wire r4_934;
assign r4_934 = in[3]? r3_1868 : r3_1867;
wire r4_935;
assign r4_935 = in[3]? r3_1870 : r3_1869;
wire r4_936;
assign r4_936 = in[3]? r3_1872 : r3_1871;
wire r4_937;
assign r4_937 = in[3]? r3_1874 : r3_1873;
wire r4_938;
assign r4_938 = in[3]? r3_1876 : r3_1875;
wire r4_939;
assign r4_939 = in[3]? r3_1878 : r3_1877;
wire r4_940;
assign r4_940 = in[3]? r3_1880 : r3_1879;
wire r4_941;
assign r4_941 = in[3]? r3_1882 : r3_1881;
wire r4_942;
assign r4_942 = in[3]? r3_1884 : r3_1883;
wire r4_943;
assign r4_943 = in[3]? r3_1886 : r3_1885;
wire r4_944;
assign r4_944 = in[3]? r3_1888 : r3_1887;
wire r4_945;
assign r4_945 = in[3]? r3_1890 : r3_1889;
wire r4_946;
assign r4_946 = in[3]? r3_1892 : r3_1891;
wire r4_947;
assign r4_947 = in[3]? r3_1894 : r3_1893;
wire r4_948;
assign r4_948 = in[3]? r3_1896 : r3_1895;
wire r4_949;
assign r4_949 = in[3]? r3_1898 : r3_1897;
wire r4_950;
assign r4_950 = in[3]? r3_1900 : r3_1899;
wire r4_951;
assign r4_951 = in[3]? r3_1902 : r3_1901;
wire r4_952;
assign r4_952 = in[3]? r3_1904 : r3_1903;
wire r4_953;
assign r4_953 = in[3]? r3_1906 : r3_1905;
wire r4_954;
assign r4_954 = in[3]? r3_1908 : r3_1907;
wire r4_955;
assign r4_955 = in[3]? r3_1910 : r3_1909;
wire r4_956;
assign r4_956 = in[3]? r3_1912 : r3_1911;
wire r4_957;
assign r4_957 = in[3]? r3_1914 : r3_1913;
wire r4_958;
assign r4_958 = in[3]? r3_1916 : r3_1915;
wire r4_959;
assign r4_959 = in[3]? r3_1918 : r3_1917;
wire r4_960;
assign r4_960 = in[3]? r3_1920 : r3_1919;
wire r4_961;
assign r4_961 = in[3]? r3_1922 : r3_1921;
wire r4_962;
assign r4_962 = in[3]? r3_1924 : r3_1923;
wire r4_963;
assign r4_963 = in[3]? r3_1926 : r3_1925;
wire r4_964;
assign r4_964 = in[3]? r3_1928 : r3_1927;
wire r4_965;
assign r4_965 = in[3]? r3_1930 : r3_1929;
wire r4_966;
assign r4_966 = in[3]? r3_1932 : r3_1931;
wire r4_967;
assign r4_967 = in[3]? r3_1934 : r3_1933;
wire r4_968;
assign r4_968 = in[3]? r3_1936 : r3_1935;
wire r4_969;
assign r4_969 = in[3]? r3_1938 : r3_1937;
wire r4_970;
assign r4_970 = in[3]? r3_1940 : r3_1939;
wire r4_971;
assign r4_971 = in[3]? r3_1942 : r3_1941;
wire r4_972;
assign r4_972 = in[3]? r3_1944 : r3_1943;
wire r4_973;
assign r4_973 = in[3]? r3_1946 : r3_1945;
wire r4_974;
assign r4_974 = in[3]? r3_1948 : r3_1947;
wire r4_975;
assign r4_975 = in[3]? r3_1950 : r3_1949;
wire r4_976;
assign r4_976 = in[3]? r3_1952 : r3_1951;
wire r4_977;
assign r4_977 = in[3]? r3_1954 : r3_1953;
wire r4_978;
assign r4_978 = in[3]? r3_1956 : r3_1955;
wire r4_979;
assign r4_979 = in[3]? r3_1958 : r3_1957;
wire r4_980;
assign r4_980 = in[3]? r3_1960 : r3_1959;
wire r4_981;
assign r4_981 = in[3]? r3_1962 : r3_1961;
wire r4_982;
assign r4_982 = in[3]? r3_1964 : r3_1963;
wire r4_983;
assign r4_983 = in[3]? r3_1966 : r3_1965;
wire r4_984;
assign r4_984 = in[3]? r3_1968 : r3_1967;
wire r4_985;
assign r4_985 = in[3]? r3_1970 : r3_1969;
wire r4_986;
assign r4_986 = in[3]? r3_1972 : r3_1971;
wire r4_987;
assign r4_987 = in[3]? r3_1974 : r3_1973;
wire r4_988;
assign r4_988 = in[3]? r3_1976 : r3_1975;
wire r4_989;
assign r4_989 = in[3]? r3_1978 : r3_1977;
wire r4_990;
assign r4_990 = in[3]? r3_1980 : r3_1979;
wire r4_991;
assign r4_991 = in[3]? r3_1982 : r3_1981;
wire r4_992;
assign r4_992 = in[3]? r3_1984 : r3_1983;
wire r4_993;
assign r4_993 = in[3]? r3_1986 : r3_1985;
wire r4_994;
assign r4_994 = in[3]? r3_1988 : r3_1987;
wire r4_995;
assign r4_995 = in[3]? r3_1990 : r3_1989;
wire r4_996;
assign r4_996 = in[3]? r3_1992 : r3_1991;
wire r4_997;
assign r4_997 = in[3]? r3_1994 : r3_1993;
wire r4_998;
assign r4_998 = in[3]? r3_1996 : r3_1995;
wire r4_999;
assign r4_999 = in[3]? r3_1998 : r3_1997;
wire r4_1000;
assign r4_1000 = in[3]? r3_2000 : r3_1999;
wire r4_1001;
assign r4_1001 = in[3]? r3_2002 : r3_2001;
wire r4_1002;
assign r4_1002 = in[3]? r3_2004 : r3_2003;
wire r4_1003;
assign r4_1003 = in[3]? r3_2006 : r3_2005;
wire r4_1004;
assign r4_1004 = in[3]? r3_2008 : r3_2007;
wire r4_1005;
assign r4_1005 = in[3]? r3_2010 : r3_2009;
wire r4_1006;
assign r4_1006 = in[3]? r3_2012 : r3_2011;
wire r4_1007;
assign r4_1007 = in[3]? r3_2014 : r3_2013;
wire r4_1008;
assign r4_1008 = in[3]? r3_2016 : r3_2015;
wire r4_1009;
assign r4_1009 = in[3]? r3_2018 : r3_2017;
wire r4_1010;
assign r4_1010 = in[3]? r3_2020 : r3_2019;
wire r4_1011;
assign r4_1011 = in[3]? r3_2022 : r3_2021;
wire r4_1012;
assign r4_1012 = in[3]? r3_2024 : r3_2023;
wire r4_1013;
assign r4_1013 = in[3]? r3_2026 : r3_2025;
wire r4_1014;
assign r4_1014 = in[3]? r3_2028 : r3_2027;
wire r4_1015;
assign r4_1015 = in[3]? r3_2030 : r3_2029;
wire r4_1016;
assign r4_1016 = in[3]? r3_2032 : r3_2031;
wire r4_1017;
assign r4_1017 = in[3]? r3_2034 : r3_2033;
wire r4_1018;
assign r4_1018 = in[3]? r3_2036 : r3_2035;
wire r4_1019;
assign r4_1019 = in[3]? r3_2038 : r3_2037;
wire r4_1020;
assign r4_1020 = in[3]? r3_2040 : r3_2039;
wire r4_1021;
assign r4_1021 = in[3]? r3_2042 : r3_2041;
wire r4_1022;
assign r4_1022 = in[3]? r3_2044 : r3_2043;
wire r4_1023;
assign r4_1023 = in[3]? r3_2046 : r3_2045;
wire r4_1024;
assign r4_1024 = in[3]? r3_2048 : r3_2047;
wire r4_1025;
assign r4_1025 = in[3]? r3_2050 : r3_2049;
wire r4_1026;
assign r4_1026 = in[3]? r3_2052 : r3_2051;
wire r4_1027;
assign r4_1027 = in[3]? r3_2054 : r3_2053;
wire r4_1028;
assign r4_1028 = in[3]? r3_2056 : r3_2055;
wire r4_1029;
assign r4_1029 = in[3]? r3_2058 : r3_2057;
wire r4_1030;
assign r4_1030 = in[3]? r3_2060 : r3_2059;
wire r4_1031;
assign r4_1031 = in[3]? r3_2062 : r3_2061;
wire r4_1032;
assign r4_1032 = in[3]? r3_2064 : r3_2063;
wire r4_1033;
assign r4_1033 = in[3]? r3_2066 : r3_2065;
wire r4_1034;
assign r4_1034 = in[3]? r3_2068 : r3_2067;
wire r4_1035;
assign r4_1035 = in[3]? r3_2070 : r3_2069;
wire r4_1036;
assign r4_1036 = in[3]? r3_2072 : r3_2071;
wire r4_1037;
assign r4_1037 = in[3]? r3_2074 : r3_2073;
wire r4_1038;
assign r4_1038 = in[3]? r3_2076 : r3_2075;
wire r4_1039;
assign r4_1039 = in[3]? r3_2078 : r3_2077;
wire r4_1040;
assign r4_1040 = in[3]? r3_2080 : r3_2079;
wire r4_1041;
assign r4_1041 = in[3]? r3_2082 : r3_2081;
wire r4_1042;
assign r4_1042 = in[3]? r3_2084 : r3_2083;
wire r4_1043;
assign r4_1043 = in[3]? r3_2086 : r3_2085;
wire r4_1044;
assign r4_1044 = in[3]? r3_2088 : r3_2087;
wire r4_1045;
assign r4_1045 = in[3]? r3_2090 : r3_2089;
wire r4_1046;
assign r4_1046 = in[3]? r3_2092 : r3_2091;
wire r4_1047;
assign r4_1047 = in[3]? r3_2094 : r3_2093;
wire r4_1048;
assign r4_1048 = in[3]? r3_2096 : r3_2095;
wire r4_1049;
assign r4_1049 = in[3]? r3_2098 : r3_2097;
wire r4_1050;
assign r4_1050 = in[3]? r3_2100 : r3_2099;
wire r4_1051;
assign r4_1051 = in[3]? r3_2102 : r3_2101;
wire r4_1052;
assign r4_1052 = in[3]? r3_2104 : r3_2103;
wire r4_1053;
assign r4_1053 = in[3]? r3_2106 : r3_2105;
wire r4_1054;
assign r4_1054 = in[3]? r3_2108 : r3_2107;
wire r4_1055;
assign r4_1055 = in[3]? r3_2110 : r3_2109;
wire r4_1056;
assign r4_1056 = in[3]? r3_2112 : r3_2111;
wire r4_1057;
assign r4_1057 = in[3]? r3_2114 : r3_2113;
wire r4_1058;
assign r4_1058 = in[3]? r3_2116 : r3_2115;
wire r4_1059;
assign r4_1059 = in[3]? r3_2118 : r3_2117;
wire r4_1060;
assign r4_1060 = in[3]? r3_2120 : r3_2119;
wire r4_1061;
assign r4_1061 = in[3]? r3_2122 : r3_2121;
wire r4_1062;
assign r4_1062 = in[3]? r3_2124 : r3_2123;
wire r4_1063;
assign r4_1063 = in[3]? r3_2126 : r3_2125;
wire r4_1064;
assign r4_1064 = in[3]? r3_2128 : r3_2127;
wire r4_1065;
assign r4_1065 = in[3]? r3_2130 : r3_2129;
wire r4_1066;
assign r4_1066 = in[3]? r3_2132 : r3_2131;
wire r4_1067;
assign r4_1067 = in[3]? r3_2134 : r3_2133;
wire r4_1068;
assign r4_1068 = in[3]? r3_2136 : r3_2135;
wire r4_1069;
assign r4_1069 = in[3]? r3_2138 : r3_2137;
wire r4_1070;
assign r4_1070 = in[3]? r3_2140 : r3_2139;
wire r4_1071;
assign r4_1071 = in[3]? r3_2142 : r3_2141;
wire r4_1072;
assign r4_1072 = in[3]? r3_2144 : r3_2143;
wire r4_1073;
assign r4_1073 = in[3]? r3_2146 : r3_2145;
wire r4_1074;
assign r4_1074 = in[3]? r3_2148 : r3_2147;
wire r4_1075;
assign r4_1075 = in[3]? r3_2150 : r3_2149;
wire r4_1076;
assign r4_1076 = in[3]? r3_2152 : r3_2151;
wire r4_1077;
assign r4_1077 = in[3]? r3_2154 : r3_2153;
wire r4_1078;
assign r4_1078 = in[3]? r3_2156 : r3_2155;
wire r4_1079;
assign r4_1079 = in[3]? r3_2158 : r3_2157;
wire r4_1080;
assign r4_1080 = in[3]? r3_2160 : r3_2159;
wire r4_1081;
assign r4_1081 = in[3]? r3_2162 : r3_2161;
wire r4_1082;
assign r4_1082 = in[3]? r3_2164 : r3_2163;
wire r4_1083;
assign r4_1083 = in[3]? r3_2166 : r3_2165;
wire r4_1084;
assign r4_1084 = in[3]? r3_2168 : r3_2167;
wire r4_1085;
assign r4_1085 = in[3]? r3_2170 : r3_2169;
wire r4_1086;
assign r4_1086 = in[3]? r3_2172 : r3_2171;
wire r4_1087;
assign r4_1087 = in[3]? r3_2174 : r3_2173;
wire r4_1088;
assign r4_1088 = in[3]? r3_2176 : r3_2175;
wire r4_1089;
assign r4_1089 = in[3]? r3_2178 : r3_2177;
wire r4_1090;
assign r4_1090 = in[3]? r3_2180 : r3_2179;
wire r4_1091;
assign r4_1091 = in[3]? r3_2182 : r3_2181;
wire r4_1092;
assign r4_1092 = in[3]? r3_2184 : r3_2183;
wire r4_1093;
assign r4_1093 = in[3]? r3_2186 : r3_2185;
wire r4_1094;
assign r4_1094 = in[3]? r3_2188 : r3_2187;
wire r4_1095;
assign r4_1095 = in[3]? r3_2190 : r3_2189;
wire r4_1096;
assign r4_1096 = in[3]? r3_2192 : r3_2191;
wire r4_1097;
assign r4_1097 = in[3]? r3_2194 : r3_2193;
wire r4_1098;
assign r4_1098 = in[3]? r3_2196 : r3_2195;
wire r4_1099;
assign r4_1099 = in[3]? r3_2198 : r3_2197;
wire r4_1100;
assign r4_1100 = in[3]? r3_2200 : r3_2199;
wire r4_1101;
assign r4_1101 = in[3]? r3_2202 : r3_2201;
wire r4_1102;
assign r4_1102 = in[3]? r3_2204 : r3_2203;
wire r4_1103;
assign r4_1103 = in[3]? r3_2206 : r3_2205;
wire r4_1104;
assign r4_1104 = in[3]? r3_2208 : r3_2207;
wire r4_1105;
assign r4_1105 = in[3]? r3_2210 : r3_2209;
wire r4_1106;
assign r4_1106 = in[3]? r3_2212 : r3_2211;
wire r4_1107;
assign r4_1107 = in[3]? r3_2214 : r3_2213;
wire r4_1108;
assign r4_1108 = in[3]? r3_2216 : r3_2215;
wire r4_1109;
assign r4_1109 = in[3]? r3_2218 : r3_2217;
wire r4_1110;
assign r4_1110 = in[3]? r3_2220 : r3_2219;
wire r4_1111;
assign r4_1111 = in[3]? r3_2222 : r3_2221;
wire r4_1112;
assign r4_1112 = in[3]? r3_2224 : r3_2223;
wire r4_1113;
assign r4_1113 = in[3]? r3_2226 : r3_2225;
wire r4_1114;
assign r4_1114 = in[3]? r3_2228 : r3_2227;
wire r4_1115;
assign r4_1115 = in[3]? r3_2230 : r3_2229;
wire r4_1116;
assign r4_1116 = in[3]? r3_2232 : r3_2231;
wire r4_1117;
assign r4_1117 = in[3]? r3_2234 : r3_2233;
wire r4_1118;
assign r4_1118 = in[3]? r3_2236 : r3_2235;
wire r4_1119;
assign r4_1119 = in[3]? r3_2238 : r3_2237;
wire r4_1120;
assign r4_1120 = in[3]? r3_2240 : r3_2239;
wire r4_1121;
assign r4_1121 = in[3]? r3_2242 : r3_2241;
wire r4_1122;
assign r4_1122 = in[3]? r3_2244 : r3_2243;
wire r4_1123;
assign r4_1123 = in[3]? r3_2246 : r3_2245;
wire r4_1124;
assign r4_1124 = in[3]? r3_2248 : r3_2247;
wire r4_1125;
assign r4_1125 = in[3]? r3_2250 : r3_2249;
wire r4_1126;
assign r4_1126 = in[3]? r3_2252 : r3_2251;
wire r4_1127;
assign r4_1127 = in[3]? r3_2254 : r3_2253;
wire r4_1128;
assign r4_1128 = in[3]? r3_2256 : r3_2255;
wire r4_1129;
assign r4_1129 = in[3]? r3_2258 : r3_2257;
wire r4_1130;
assign r4_1130 = in[3]? r3_2260 : r3_2259;
wire r4_1131;
assign r4_1131 = in[3]? r3_2262 : r3_2261;
wire r4_1132;
assign r4_1132 = in[3]? r3_2264 : r3_2263;
wire r4_1133;
assign r4_1133 = in[3]? r3_2266 : r3_2265;
wire r4_1134;
assign r4_1134 = in[3]? r3_2268 : r3_2267;
wire r4_1135;
assign r4_1135 = in[3]? r3_2270 : r3_2269;
wire r4_1136;
assign r4_1136 = in[3]? r3_2272 : r3_2271;
wire r4_1137;
assign r4_1137 = in[3]? r3_2274 : r3_2273;
wire r4_1138;
assign r4_1138 = in[3]? r3_2276 : r3_2275;
wire r4_1139;
assign r4_1139 = in[3]? r3_2278 : r3_2277;
wire r4_1140;
assign r4_1140 = in[3]? r3_2280 : r3_2279;
wire r4_1141;
assign r4_1141 = in[3]? r3_2282 : r3_2281;
wire r4_1142;
assign r4_1142 = in[3]? r3_2284 : r3_2283;
wire r4_1143;
assign r4_1143 = in[3]? r3_2286 : r3_2285;
wire r4_1144;
assign r4_1144 = in[3]? r3_2288 : r3_2287;
wire r4_1145;
assign r4_1145 = in[3]? r3_2290 : r3_2289;
wire r4_1146;
assign r4_1146 = in[3]? r3_2292 : r3_2291;
wire r4_1147;
assign r4_1147 = in[3]? r3_2294 : r3_2293;
wire r4_1148;
assign r4_1148 = in[3]? r3_2296 : r3_2295;
wire r4_1149;
assign r4_1149 = in[3]? r3_2298 : r3_2297;
wire r4_1150;
assign r4_1150 = in[3]? r3_2300 : r3_2299;
wire r4_1151;
assign r4_1151 = in[3]? r3_2302 : r3_2301;
wire r4_1152;
assign r4_1152 = in[3]? r3_2304 : r3_2303;
wire r4_1153;
assign r4_1153 = in[3]? r3_2306 : r3_2305;
wire r4_1154;
assign r4_1154 = in[3]? r3_2308 : r3_2307;
wire r4_1155;
assign r4_1155 = in[3]? r3_2310 : r3_2309;
wire r4_1156;
assign r4_1156 = in[3]? r3_2312 : r3_2311;
wire r4_1157;
assign r4_1157 = in[3]? r3_2314 : r3_2313;
wire r4_1158;
assign r4_1158 = in[3]? r3_2316 : r3_2315;
wire r4_1159;
assign r4_1159 = in[3]? r3_2318 : r3_2317;
wire r4_1160;
assign r4_1160 = in[3]? r3_2320 : r3_2319;
wire r4_1161;
assign r4_1161 = in[3]? r3_2322 : r3_2321;
wire r4_1162;
assign r4_1162 = in[3]? r3_2324 : r3_2323;
wire r4_1163;
assign r4_1163 = in[3]? r3_2326 : r3_2325;
wire r4_1164;
assign r4_1164 = in[3]? r3_2328 : r3_2327;
wire r4_1165;
assign r4_1165 = in[3]? r3_2330 : r3_2329;
wire r4_1166;
assign r4_1166 = in[3]? r3_2332 : r3_2331;
wire r4_1167;
assign r4_1167 = in[3]? r3_2334 : r3_2333;
wire r4_1168;
assign r4_1168 = in[3]? r3_2336 : r3_2335;
wire r4_1169;
assign r4_1169 = in[3]? r3_2338 : r3_2337;
wire r4_1170;
assign r4_1170 = in[3]? r3_2340 : r3_2339;
wire r4_1171;
assign r4_1171 = in[3]? r3_2342 : r3_2341;
wire r4_1172;
assign r4_1172 = in[3]? r3_2344 : r3_2343;
wire r4_1173;
assign r4_1173 = in[3]? r3_2346 : r3_2345;
wire r4_1174;
assign r4_1174 = in[3]? r3_2348 : r3_2347;
wire r4_1175;
assign r4_1175 = in[3]? r3_2350 : r3_2349;
wire r4_1176;
assign r4_1176 = in[3]? r3_2352 : r3_2351;
wire r4_1177;
assign r4_1177 = in[3]? r3_2354 : r3_2353;
wire r4_1178;
assign r4_1178 = in[3]? r3_2356 : r3_2355;
wire r4_1179;
assign r4_1179 = in[3]? r3_2358 : r3_2357;
wire r4_1180;
assign r4_1180 = in[3]? r3_2360 : r3_2359;
wire r4_1181;
assign r4_1181 = in[3]? r3_2362 : r3_2361;
wire r4_1182;
assign r4_1182 = in[3]? r3_2364 : r3_2363;
wire r4_1183;
assign r4_1183 = in[3]? r3_2366 : r3_2365;
wire r4_1184;
assign r4_1184 = in[3]? r3_2368 : r3_2367;
wire r4_1185;
assign r4_1185 = in[3]? r3_2370 : r3_2369;
wire r4_1186;
assign r4_1186 = in[3]? r3_2372 : r3_2371;
wire r4_1187;
assign r4_1187 = in[3]? r3_2374 : r3_2373;
wire r4_1188;
assign r4_1188 = in[3]? r3_2376 : r3_2375;
wire r4_1189;
assign r4_1189 = in[3]? r3_2378 : r3_2377;
wire r4_1190;
assign r4_1190 = in[3]? r3_2380 : r3_2379;
wire r4_1191;
assign r4_1191 = in[3]? r3_2382 : r3_2381;
wire r4_1192;
assign r4_1192 = in[3]? r3_2384 : r3_2383;
wire r4_1193;
assign r4_1193 = in[3]? r3_2386 : r3_2385;
wire r4_1194;
assign r4_1194 = in[3]? r3_2388 : r3_2387;
wire r4_1195;
assign r4_1195 = in[3]? r3_2390 : r3_2389;
wire r4_1196;
assign r4_1196 = in[3]? r3_2392 : r3_2391;
wire r4_1197;
assign r4_1197 = in[3]? r3_2394 : r3_2393;
wire r4_1198;
assign r4_1198 = in[3]? r3_2396 : r3_2395;
wire r4_1199;
assign r4_1199 = in[3]? r3_2398 : r3_2397;
wire r4_1200;
assign r4_1200 = in[3]? r3_2400 : r3_2399;
wire r4_1201;
assign r4_1201 = in[3]? r3_2402 : r3_2401;
wire r4_1202;
assign r4_1202 = in[3]? r3_2404 : r3_2403;
wire r4_1203;
assign r4_1203 = in[3]? r3_2406 : r3_2405;
wire r4_1204;
assign r4_1204 = in[3]? r3_2408 : r3_2407;
wire r4_1205;
assign r4_1205 = in[3]? r3_2410 : r3_2409;
wire r4_1206;
assign r4_1206 = in[3]? r3_2412 : r3_2411;
wire r4_1207;
assign r4_1207 = in[3]? r3_2414 : r3_2413;
wire r4_1208;
assign r4_1208 = in[3]? r3_2416 : r3_2415;
wire r4_1209;
assign r4_1209 = in[3]? r3_2418 : r3_2417;
wire r4_1210;
assign r4_1210 = in[3]? r3_2420 : r3_2419;
wire r4_1211;
assign r4_1211 = in[3]? r3_2422 : r3_2421;
wire r4_1212;
assign r4_1212 = in[3]? r3_2424 : r3_2423;
wire r4_1213;
assign r4_1213 = in[3]? r3_2426 : r3_2425;
wire r4_1214;
assign r4_1214 = in[3]? r3_2428 : r3_2427;
wire r4_1215;
assign r4_1215 = in[3]? r3_2430 : r3_2429;
wire r4_1216;
assign r4_1216 = in[3]? r3_2432 : r3_2431;
wire r4_1217;
assign r4_1217 = in[3]? r3_2434 : r3_2433;
wire r4_1218;
assign r4_1218 = in[3]? r3_2436 : r3_2435;
wire r4_1219;
assign r4_1219 = in[3]? r3_2438 : r3_2437;
wire r4_1220;
assign r4_1220 = in[3]? r3_2440 : r3_2439;
wire r4_1221;
assign r4_1221 = in[3]? r3_2442 : r3_2441;
wire r4_1222;
assign r4_1222 = in[3]? r3_2444 : r3_2443;
wire r4_1223;
assign r4_1223 = in[3]? r3_2446 : r3_2445;
wire r4_1224;
assign r4_1224 = in[3]? r3_2448 : r3_2447;
wire r4_1225;
assign r4_1225 = in[3]? r3_2450 : r3_2449;
wire r4_1226;
assign r4_1226 = in[3]? r3_2452 : r3_2451;
wire r4_1227;
assign r4_1227 = in[3]? r3_2454 : r3_2453;
wire r4_1228;
assign r4_1228 = in[3]? r3_2456 : r3_2455;
wire r4_1229;
assign r4_1229 = in[3]? r3_2458 : r3_2457;
wire r4_1230;
assign r4_1230 = in[3]? r3_2460 : r3_2459;
wire r4_1231;
assign r4_1231 = in[3]? r3_2462 : r3_2461;
wire r4_1232;
assign r4_1232 = in[3]? r3_2464 : r3_2463;
wire r4_1233;
assign r4_1233 = in[3]? r3_2466 : r3_2465;
wire r4_1234;
assign r4_1234 = in[3]? r3_2468 : r3_2467;
wire r4_1235;
assign r4_1235 = in[3]? r3_2470 : r3_2469;
wire r4_1236;
assign r4_1236 = in[3]? r3_2472 : r3_2471;
wire r4_1237;
assign r4_1237 = in[3]? r3_2474 : r3_2473;
wire r4_1238;
assign r4_1238 = in[3]? r3_2476 : r3_2475;
wire r4_1239;
assign r4_1239 = in[3]? r3_2478 : r3_2477;
wire r4_1240;
assign r4_1240 = in[3]? r3_2480 : r3_2479;
wire r4_1241;
assign r4_1241 = in[3]? r3_2482 : r3_2481;
wire r4_1242;
assign r4_1242 = in[3]? r3_2484 : r3_2483;
wire r4_1243;
assign r4_1243 = in[3]? r3_2486 : r3_2485;
wire r4_1244;
assign r4_1244 = in[3]? r3_2488 : r3_2487;
wire r4_1245;
assign r4_1245 = in[3]? r3_2490 : r3_2489;
wire r4_1246;
assign r4_1246 = in[3]? r3_2492 : r3_2491;
wire r4_1247;
assign r4_1247 = in[3]? r3_2494 : r3_2493;
wire r4_1248;
assign r4_1248 = in[3]? r3_2496 : r3_2495;
wire r4_1249;
assign r4_1249 = in[3]? r3_2498 : r3_2497;
wire r4_1250;
assign r4_1250 = in[3]? r3_2500 : r3_2499;
wire r4_1251;
assign r4_1251 = in[3]? r3_2502 : r3_2501;
wire r4_1252;
assign r4_1252 = in[3]? r3_2504 : r3_2503;
wire r4_1253;
assign r4_1253 = in[3]? r3_2506 : r3_2505;
wire r4_1254;
assign r4_1254 = in[3]? r3_2508 : r3_2507;
wire r4_1255;
assign r4_1255 = in[3]? r3_2510 : r3_2509;
wire r4_1256;
assign r4_1256 = in[3]? r3_2512 : r3_2511;
wire r4_1257;
assign r4_1257 = in[3]? r3_2514 : r3_2513;
wire r4_1258;
assign r4_1258 = in[3]? r3_2516 : r3_2515;
wire r4_1259;
assign r4_1259 = in[3]? r3_2518 : r3_2517;
wire r4_1260;
assign r4_1260 = in[3]? r3_2520 : r3_2519;
wire r4_1261;
assign r4_1261 = in[3]? r3_2522 : r3_2521;
wire r4_1262;
assign r4_1262 = in[3]? r3_2524 : r3_2523;
wire r4_1263;
assign r4_1263 = in[3]? r3_2526 : r3_2525;
wire r4_1264;
assign r4_1264 = in[3]? r3_2528 : r3_2527;
wire r4_1265;
assign r4_1265 = in[3]? r3_2530 : r3_2529;
wire r4_1266;
assign r4_1266 = in[3]? r3_2532 : r3_2531;
wire r4_1267;
assign r4_1267 = in[3]? r3_2534 : r3_2533;
wire r4_1268;
assign r4_1268 = in[3]? r3_2536 : r3_2535;
wire r4_1269;
assign r4_1269 = in[3]? r3_2538 : r3_2537;
wire r4_1270;
assign r4_1270 = in[3]? r3_2540 : r3_2539;
wire r4_1271;
assign r4_1271 = in[3]? r3_2542 : r3_2541;
wire r4_1272;
assign r4_1272 = in[3]? r3_2544 : r3_2543;
wire r4_1273;
assign r4_1273 = in[3]? r3_2546 : r3_2545;
wire r4_1274;
assign r4_1274 = in[3]? r3_2548 : r3_2547;
wire r4_1275;
assign r4_1275 = in[3]? r3_2550 : r3_2549;
wire r4_1276;
assign r4_1276 = in[3]? r3_2552 : r3_2551;
wire r4_1277;
assign r4_1277 = in[3]? r3_2554 : r3_2553;
wire r4_1278;
assign r4_1278 = in[3]? r3_2556 : r3_2555;
wire r4_1279;
assign r4_1279 = in[3]? r3_2558 : r3_2557;
wire r4_1280;
assign r4_1280 = in[3]? r3_2560 : r3_2559;
wire r4_1281;
assign r4_1281 = in[3]? r3_2562 : r3_2561;
wire r4_1282;
assign r4_1282 = in[3]? r3_2564 : r3_2563;
wire r4_1283;
assign r4_1283 = in[3]? r3_2566 : r3_2565;
wire r4_1284;
assign r4_1284 = in[3]? r3_2568 : r3_2567;
wire r5_1;
assign r5_1 = in[4]? r4_2 : r4_1;
wire r5_2;
assign r5_2 = in[4]? r4_4 : r4_3;
wire r5_3;
assign r5_3 = in[4]? r4_6 : r4_5;
wire r5_4;
assign r5_4 = in[4]? r4_8 : r4_7;
wire r5_5;
assign r5_5 = in[4]? r4_10 : r4_9;
wire r5_6;
assign r5_6 = in[4]? r4_12 : r4_11;
wire r5_7;
assign r5_7 = in[4]? r4_14 : r4_13;
wire r5_8;
assign r5_8 = in[4]? r4_16 : r4_15;
wire r5_9;
assign r5_9 = in[4]? r4_18 : r4_17;
wire r5_10;
assign r5_10 = in[4]? r4_20 : r4_19;
wire r5_11;
assign r5_11 = in[4]? r4_22 : r4_21;
wire r5_12;
assign r5_12 = in[4]? r4_24 : r4_23;
wire r5_13;
assign r5_13 = in[4]? r4_26 : r4_25;
wire r5_14;
assign r5_14 = in[4]? r4_28 : r4_27;
wire r5_15;
assign r5_15 = in[4]? r4_30 : r4_29;
wire r5_16;
assign r5_16 = in[4]? r4_32 : r4_31;
wire r5_17;
assign r5_17 = in[4]? r4_34 : r4_33;
wire r5_18;
assign r5_18 = in[4]? r4_36 : r4_35;
wire r5_19;
assign r5_19 = in[4]? r4_38 : r4_37;
wire r5_20;
assign r5_20 = in[4]? r4_40 : r4_39;
wire r5_21;
assign r5_21 = in[4]? r4_42 : r4_41;
wire r5_22;
assign r5_22 = in[4]? r4_44 : r4_43;
wire r5_23;
assign r5_23 = in[4]? r4_46 : r4_45;
wire r5_24;
assign r5_24 = in[4]? r4_48 : r4_47;
wire r5_25;
assign r5_25 = in[4]? r4_50 : r4_49;
wire r5_26;
assign r5_26 = in[4]? r4_52 : r4_51;
wire r5_27;
assign r5_27 = in[4]? r4_54 : r4_53;
wire r5_28;
assign r5_28 = in[4]? r4_56 : r4_55;
wire r5_29;
assign r5_29 = in[4]? r4_58 : r4_57;
wire r5_30;
assign r5_30 = in[4]? r4_60 : r4_59;
wire r5_31;
assign r5_31 = in[4]? r4_62 : r4_61;
wire r5_32;
assign r5_32 = in[4]? r4_64 : r4_63;
wire r5_33;
assign r5_33 = in[4]? r4_66 : r4_65;
wire r5_34;
assign r5_34 = in[4]? r4_68 : r4_67;
wire r5_35;
assign r5_35 = in[4]? r4_70 : r4_69;
wire r5_36;
assign r5_36 = in[4]? r4_72 : r4_71;
wire r5_37;
assign r5_37 = in[4]? r4_74 : r4_73;
wire r5_38;
assign r5_38 = in[4]? r4_76 : r4_75;
wire r5_39;
assign r5_39 = in[4]? r4_78 : r4_77;
wire r5_40;
assign r5_40 = in[4]? r4_80 : r4_79;
wire r5_41;
assign r5_41 = in[4]? r4_82 : r4_81;
wire r5_42;
assign r5_42 = in[4]? r4_84 : r4_83;
wire r5_43;
assign r5_43 = in[4]? r4_86 : r4_85;
wire r5_44;
assign r5_44 = in[4]? r4_88 : r4_87;
wire r5_45;
assign r5_45 = in[4]? r4_90 : r4_89;
wire r5_46;
assign r5_46 = in[4]? r4_92 : r4_91;
wire r5_47;
assign r5_47 = in[4]? r4_94 : r4_93;
wire r5_48;
assign r5_48 = in[4]? r4_96 : r4_95;
wire r5_49;
assign r5_49 = in[4]? r4_98 : r4_97;
wire r5_50;
assign r5_50 = in[4]? r4_100 : r4_99;
wire r5_51;
assign r5_51 = in[4]? r4_102 : r4_101;
wire r5_52;
assign r5_52 = in[4]? r4_104 : r4_103;
wire r5_53;
assign r5_53 = in[4]? r4_106 : r4_105;
wire r5_54;
assign r5_54 = in[4]? r4_108 : r4_107;
wire r5_55;
assign r5_55 = in[4]? r4_110 : r4_109;
wire r5_56;
assign r5_56 = in[4]? r4_112 : r4_111;
wire r5_57;
assign r5_57 = in[4]? r4_114 : r4_113;
wire r5_58;
assign r5_58 = in[4]? r4_116 : r4_115;
wire r5_59;
assign r5_59 = in[4]? r4_118 : r4_117;
wire r5_60;
assign r5_60 = in[4]? r4_120 : r4_119;
wire r5_61;
assign r5_61 = in[4]? r4_122 : r4_121;
wire r5_62;
assign r5_62 = in[4]? r4_124 : r4_123;
wire r5_63;
assign r5_63 = in[4]? r4_126 : r4_125;
wire r5_64;
assign r5_64 = in[4]? r4_128 : r4_127;
wire r5_65;
assign r5_65 = in[4]? r4_130 : r4_129;
wire r5_66;
assign r5_66 = in[4]? r4_132 : r4_131;
wire r5_67;
assign r5_67 = in[4]? r4_134 : r4_133;
wire r5_68;
assign r5_68 = in[4]? r4_136 : r4_135;
wire r5_69;
assign r5_69 = in[4]? r4_138 : r4_137;
wire r5_70;
assign r5_70 = in[4]? r4_140 : r4_139;
wire r5_71;
assign r5_71 = in[4]? r4_142 : r4_141;
wire r5_72;
assign r5_72 = in[4]? r4_144 : r4_143;
wire r5_73;
assign r5_73 = in[4]? r4_146 : r4_145;
wire r5_74;
assign r5_74 = in[4]? r4_148 : r4_147;
wire r5_75;
assign r5_75 = in[4]? r4_150 : r4_149;
wire r5_76;
assign r5_76 = in[4]? r4_152 : r4_151;
wire r5_77;
assign r5_77 = in[4]? r4_154 : r4_153;
wire r5_78;
assign r5_78 = in[4]? r4_156 : r4_155;
wire r5_79;
assign r5_79 = in[4]? r4_158 : r4_157;
wire r5_80;
assign r5_80 = in[4]? r4_160 : r4_159;
wire r5_81;
assign r5_81 = in[4]? r4_162 : r4_161;
wire r5_82;
assign r5_82 = in[4]? r4_164 : r4_163;
wire r5_83;
assign r5_83 = in[4]? r4_166 : r4_165;
wire r5_84;
assign r5_84 = in[4]? r4_168 : r4_167;
wire r5_85;
assign r5_85 = in[4]? r4_170 : r4_169;
wire r5_86;
assign r5_86 = in[4]? r4_172 : r4_171;
wire r5_87;
assign r5_87 = in[4]? r4_174 : r4_173;
wire r5_88;
assign r5_88 = in[4]? r4_176 : r4_175;
wire r5_89;
assign r5_89 = in[4]? r4_178 : r4_177;
wire r5_90;
assign r5_90 = in[4]? r4_180 : r4_179;
wire r5_91;
assign r5_91 = in[4]? r4_182 : r4_181;
wire r5_92;
assign r5_92 = in[4]? r4_184 : r4_183;
wire r5_93;
assign r5_93 = in[4]? r4_186 : r4_185;
wire r5_94;
assign r5_94 = in[4]? r4_188 : r4_187;
wire r5_95;
assign r5_95 = in[4]? r4_190 : r4_189;
wire r5_96;
assign r5_96 = in[4]? r4_192 : r4_191;
wire r5_97;
assign r5_97 = in[4]? r4_194 : r4_193;
wire r5_98;
assign r5_98 = in[4]? r4_196 : r4_195;
wire r5_99;
assign r5_99 = in[4]? r4_198 : r4_197;
wire r5_100;
assign r5_100 = in[4]? r4_200 : r4_199;
wire r5_101;
assign r5_101 = in[4]? r4_202 : r4_201;
wire r5_102;
assign r5_102 = in[4]? r4_204 : r4_203;
wire r5_103;
assign r5_103 = in[4]? r4_206 : r4_205;
wire r5_104;
assign r5_104 = in[4]? r4_208 : r4_207;
wire r5_105;
assign r5_105 = in[4]? r4_210 : r4_209;
wire r5_106;
assign r5_106 = in[4]? r4_212 : r4_211;
wire r5_107;
assign r5_107 = in[4]? r4_214 : r4_213;
wire r5_108;
assign r5_108 = in[4]? r4_216 : r4_215;
wire r5_109;
assign r5_109 = in[4]? r4_218 : r4_217;
wire r5_110;
assign r5_110 = in[4]? r4_220 : r4_219;
wire r5_111;
assign r5_111 = in[4]? r4_222 : r4_221;
wire r5_112;
assign r5_112 = in[4]? r4_224 : r4_223;
wire r5_113;
assign r5_113 = in[4]? r4_226 : r4_225;
wire r5_114;
assign r5_114 = in[4]? r4_228 : r4_227;
wire r5_115;
assign r5_115 = in[4]? r4_230 : r4_229;
wire r5_116;
assign r5_116 = in[4]? r4_232 : r4_231;
wire r5_117;
assign r5_117 = in[4]? r4_234 : r4_233;
wire r5_118;
assign r5_118 = in[4]? r4_236 : r4_235;
wire r5_119;
assign r5_119 = in[4]? r4_238 : r4_237;
wire r5_120;
assign r5_120 = in[4]? r4_240 : r4_239;
wire r5_121;
assign r5_121 = in[4]? r4_242 : r4_241;
wire r5_122;
assign r5_122 = in[4]? r4_244 : r4_243;
wire r5_123;
assign r5_123 = in[4]? r4_246 : r4_245;
wire r5_124;
assign r5_124 = in[4]? r4_248 : r4_247;
wire r5_125;
assign r5_125 = in[4]? r4_250 : r4_249;
wire r5_126;
assign r5_126 = in[4]? r4_252 : r4_251;
wire r5_127;
assign r5_127 = in[4]? r4_254 : r4_253;
wire r5_128;
assign r5_128 = in[4]? r4_256 : r4_255;
wire r5_129;
assign r5_129 = in[4]? r4_258 : r4_257;
wire r5_130;
assign r5_130 = in[4]? r4_260 : r4_259;
wire r5_131;
assign r5_131 = in[4]? r4_262 : r4_261;
wire r5_132;
assign r5_132 = in[4]? r4_264 : r4_263;
wire r5_133;
assign r5_133 = in[4]? r4_266 : r4_265;
wire r5_134;
assign r5_134 = in[4]? r4_268 : r4_267;
wire r5_135;
assign r5_135 = in[4]? r4_270 : r4_269;
wire r5_136;
assign r5_136 = in[4]? r4_272 : r4_271;
wire r5_137;
assign r5_137 = in[4]? r4_274 : r4_273;
wire r5_138;
assign r5_138 = in[4]? r4_276 : r4_275;
wire r5_139;
assign r5_139 = in[4]? r4_278 : r4_277;
wire r5_140;
assign r5_140 = in[4]? r4_280 : r4_279;
wire r5_141;
assign r5_141 = in[4]? r4_282 : r4_281;
wire r5_142;
assign r5_142 = in[4]? r4_284 : r4_283;
wire r5_143;
assign r5_143 = in[4]? r4_286 : r4_285;
wire r5_144;
assign r5_144 = in[4]? r4_288 : r4_287;
wire r5_145;
assign r5_145 = in[4]? r4_290 : r4_289;
wire r5_146;
assign r5_146 = in[4]? r4_292 : r4_291;
wire r5_147;
assign r5_147 = in[4]? r4_294 : r4_293;
wire r5_148;
assign r5_148 = in[4]? r4_296 : r4_295;
wire r5_149;
assign r5_149 = in[4]? r4_298 : r4_297;
wire r5_150;
assign r5_150 = in[4]? r4_300 : r4_299;
wire r5_151;
assign r5_151 = in[4]? r4_302 : r4_301;
wire r5_152;
assign r5_152 = in[4]? r4_304 : r4_303;
wire r5_153;
assign r5_153 = in[4]? r4_306 : r4_305;
wire r5_154;
assign r5_154 = in[4]? r4_308 : r4_307;
wire r5_155;
assign r5_155 = in[4]? r4_310 : r4_309;
wire r5_156;
assign r5_156 = in[4]? r4_312 : r4_311;
wire r5_157;
assign r5_157 = in[4]? r4_314 : r4_313;
wire r5_158;
assign r5_158 = in[4]? r4_316 : r4_315;
wire r5_159;
assign r5_159 = in[4]? r4_318 : r4_317;
wire r5_160;
assign r5_160 = in[4]? r4_320 : r4_319;
wire r5_161;
assign r5_161 = in[4]? r4_322 : r4_321;
wire r5_162;
assign r5_162 = in[4]? r4_324 : r4_323;
wire r5_163;
assign r5_163 = in[4]? r4_326 : r4_325;
wire r5_164;
assign r5_164 = in[4]? r4_328 : r4_327;
wire r5_165;
assign r5_165 = in[4]? r4_330 : r4_329;
wire r5_166;
assign r5_166 = in[4]? r4_332 : r4_331;
wire r5_167;
assign r5_167 = in[4]? r4_334 : r4_333;
wire r5_168;
assign r5_168 = in[4]? r4_336 : r4_335;
wire r5_169;
assign r5_169 = in[4]? r4_338 : r4_337;
wire r5_170;
assign r5_170 = in[4]? r4_340 : r4_339;
wire r5_171;
assign r5_171 = in[4]? r4_342 : r4_341;
wire r5_172;
assign r5_172 = in[4]? r4_344 : r4_343;
wire r5_173;
assign r5_173 = in[4]? r4_346 : r4_345;
wire r5_174;
assign r5_174 = in[4]? r4_348 : r4_347;
wire r5_175;
assign r5_175 = in[4]? r4_350 : r4_349;
wire r5_176;
assign r5_176 = in[4]? r4_352 : r4_351;
wire r5_177;
assign r5_177 = in[4]? r4_354 : r4_353;
wire r5_178;
assign r5_178 = in[4]? r4_356 : r4_355;
wire r5_179;
assign r5_179 = in[4]? r4_358 : r4_357;
wire r5_180;
assign r5_180 = in[4]? r4_360 : r4_359;
wire r5_181;
assign r5_181 = in[4]? r4_362 : r4_361;
wire r5_182;
assign r5_182 = in[4]? r4_364 : r4_363;
wire r5_183;
assign r5_183 = in[4]? r4_366 : r4_365;
wire r5_184;
assign r5_184 = in[4]? r4_368 : r4_367;
wire r5_185;
assign r5_185 = in[4]? r4_370 : r4_369;
wire r5_186;
assign r5_186 = in[4]? r4_372 : r4_371;
wire r5_187;
assign r5_187 = in[4]? r4_374 : r4_373;
wire r5_188;
assign r5_188 = in[4]? r4_376 : r4_375;
wire r5_189;
assign r5_189 = in[4]? r4_378 : r4_377;
wire r5_190;
assign r5_190 = in[4]? r4_380 : r4_379;
wire r5_191;
assign r5_191 = in[4]? r4_382 : r4_381;
wire r5_192;
assign r5_192 = in[4]? r4_384 : r4_383;
wire r5_193;
assign r5_193 = in[4]? r4_386 : r4_385;
wire r5_194;
assign r5_194 = in[4]? r4_388 : r4_387;
wire r5_195;
assign r5_195 = in[4]? r4_390 : r4_389;
wire r5_196;
assign r5_196 = in[4]? r4_392 : r4_391;
wire r5_197;
assign r5_197 = in[4]? r4_394 : r4_393;
wire r5_198;
assign r5_198 = in[4]? r4_396 : r4_395;
wire r5_199;
assign r5_199 = in[4]? r4_398 : r4_397;
wire r5_200;
assign r5_200 = in[4]? r4_400 : r4_399;
wire r5_201;
assign r5_201 = in[4]? r4_402 : r4_401;
wire r5_202;
assign r5_202 = in[4]? r4_404 : r4_403;
wire r5_203;
assign r5_203 = in[4]? r4_406 : r4_405;
wire r5_204;
assign r5_204 = in[4]? r4_408 : r4_407;
wire r5_205;
assign r5_205 = in[4]? r4_410 : r4_409;
wire r5_206;
assign r5_206 = in[4]? r4_412 : r4_411;
wire r5_207;
assign r5_207 = in[4]? r4_414 : r4_413;
wire r5_208;
assign r5_208 = in[4]? r4_416 : r4_415;
wire r5_209;
assign r5_209 = in[4]? r4_418 : r4_417;
wire r5_210;
assign r5_210 = in[4]? r4_420 : r4_419;
wire r5_211;
assign r5_211 = in[4]? r4_422 : r4_421;
wire r5_212;
assign r5_212 = in[4]? r4_424 : r4_423;
wire r5_213;
assign r5_213 = in[4]? r4_426 : r4_425;
wire r5_214;
assign r5_214 = in[4]? r4_428 : r4_427;
wire r5_215;
assign r5_215 = in[4]? r4_430 : r4_429;
wire r5_216;
assign r5_216 = in[4]? r4_432 : r4_431;
wire r5_217;
assign r5_217 = in[4]? r4_434 : r4_433;
wire r5_218;
assign r5_218 = in[4]? r4_436 : r4_435;
wire r5_219;
assign r5_219 = in[4]? r4_438 : r4_437;
wire r5_220;
assign r5_220 = in[4]? r4_440 : r4_439;
wire r5_221;
assign r5_221 = in[4]? r4_442 : r4_441;
wire r5_222;
assign r5_222 = in[4]? r4_444 : r4_443;
wire r5_223;
assign r5_223 = in[4]? r4_446 : r4_445;
wire r5_224;
assign r5_224 = in[4]? r4_448 : r4_447;
wire r5_225;
assign r5_225 = in[4]? r4_450 : r4_449;
wire r5_226;
assign r5_226 = in[4]? r4_452 : r4_451;
wire r5_227;
assign r5_227 = in[4]? r4_454 : r4_453;
wire r5_228;
assign r5_228 = in[4]? r4_456 : r4_455;
wire r5_229;
assign r5_229 = in[4]? r4_458 : r4_457;
wire r5_230;
assign r5_230 = in[4]? r4_460 : r4_459;
wire r5_231;
assign r5_231 = in[4]? r4_462 : r4_461;
wire r5_232;
assign r5_232 = in[4]? r4_464 : r4_463;
wire r5_233;
assign r5_233 = in[4]? r4_466 : r4_465;
wire r5_234;
assign r5_234 = in[4]? r4_468 : r4_467;
wire r5_235;
assign r5_235 = in[4]? r4_470 : r4_469;
wire r5_236;
assign r5_236 = in[4]? r4_472 : r4_471;
wire r5_237;
assign r5_237 = in[4]? r4_474 : r4_473;
wire r5_238;
assign r5_238 = in[4]? r4_476 : r4_475;
wire r5_239;
assign r5_239 = in[4]? r4_478 : r4_477;
wire r5_240;
assign r5_240 = in[4]? r4_480 : r4_479;
wire r5_241;
assign r5_241 = in[4]? r4_482 : r4_481;
wire r5_242;
assign r5_242 = in[4]? r4_484 : r4_483;
wire r5_243;
assign r5_243 = in[4]? r4_486 : r4_485;
wire r5_244;
assign r5_244 = in[4]? r4_488 : r4_487;
wire r5_245;
assign r5_245 = in[4]? r4_490 : r4_489;
wire r5_246;
assign r5_246 = in[4]? r4_492 : r4_491;
wire r5_247;
assign r5_247 = in[4]? r4_494 : r4_493;
wire r5_248;
assign r5_248 = in[4]? r4_496 : r4_495;
wire r5_249;
assign r5_249 = in[4]? r4_498 : r4_497;
wire r5_250;
assign r5_250 = in[4]? r4_500 : r4_499;
wire r5_251;
assign r5_251 = in[4]? r4_502 : r4_501;
wire r5_252;
assign r5_252 = in[4]? r4_504 : r4_503;
wire r5_253;
assign r5_253 = in[4]? r4_506 : r4_505;
wire r5_254;
assign r5_254 = in[4]? r4_508 : r4_507;
wire r5_255;
assign r5_255 = in[4]? r4_510 : r4_509;
wire r5_256;
assign r5_256 = in[4]? r4_512 : r4_511;
wire r5_257;
assign r5_257 = in[4]? r4_514 : r4_513;
wire r5_258;
assign r5_258 = in[4]? r4_516 : r4_515;
wire r5_259;
assign r5_259 = in[4]? r4_518 : r4_517;
wire r5_260;
assign r5_260 = in[4]? r4_520 : r4_519;
wire r5_261;
assign r5_261 = in[4]? r4_522 : r4_521;
wire r5_262;
assign r5_262 = in[4]? r4_524 : r4_523;
wire r5_263;
assign r5_263 = in[4]? r4_526 : r4_525;
wire r5_264;
assign r5_264 = in[4]? r4_528 : r4_527;
wire r5_265;
assign r5_265 = in[4]? r4_530 : r4_529;
wire r5_266;
assign r5_266 = in[4]? r4_532 : r4_531;
wire r5_267;
assign r5_267 = in[4]? r4_534 : r4_533;
wire r5_268;
assign r5_268 = in[4]? r4_536 : r4_535;
wire r5_269;
assign r5_269 = in[4]? r4_538 : r4_537;
wire r5_270;
assign r5_270 = in[4]? r4_540 : r4_539;
wire r5_271;
assign r5_271 = in[4]? r4_542 : r4_541;
wire r5_272;
assign r5_272 = in[4]? r4_544 : r4_543;
wire r5_273;
assign r5_273 = in[4]? r4_546 : r4_545;
wire r5_274;
assign r5_274 = in[4]? r4_548 : r4_547;
wire r5_275;
assign r5_275 = in[4]? r4_550 : r4_549;
wire r5_276;
assign r5_276 = in[4]? r4_552 : r4_551;
wire r5_277;
assign r5_277 = in[4]? r4_554 : r4_553;
wire r5_278;
assign r5_278 = in[4]? r4_556 : r4_555;
wire r5_279;
assign r5_279 = in[4]? r4_558 : r4_557;
wire r5_280;
assign r5_280 = in[4]? r4_560 : r4_559;
wire r5_281;
assign r5_281 = in[4]? r4_562 : r4_561;
wire r5_282;
assign r5_282 = in[4]? r4_564 : r4_563;
wire r5_283;
assign r5_283 = in[4]? r4_566 : r4_565;
wire r5_284;
assign r5_284 = in[4]? r4_568 : r4_567;
wire r5_285;
assign r5_285 = in[4]? r4_570 : r4_569;
wire r5_286;
assign r5_286 = in[4]? r4_572 : r4_571;
wire r5_287;
assign r5_287 = in[4]? r4_574 : r4_573;
wire r5_288;
assign r5_288 = in[4]? r4_576 : r4_575;
wire r5_289;
assign r5_289 = in[4]? r4_578 : r4_577;
wire r5_290;
assign r5_290 = in[4]? r4_580 : r4_579;
wire r5_291;
assign r5_291 = in[4]? r4_582 : r4_581;
wire r5_292;
assign r5_292 = in[4]? r4_584 : r4_583;
wire r5_293;
assign r5_293 = in[4]? r4_586 : r4_585;
wire r5_294;
assign r5_294 = in[4]? r4_588 : r4_587;
wire r5_295;
assign r5_295 = in[4]? r4_590 : r4_589;
wire r5_296;
assign r5_296 = in[4]? r4_592 : r4_591;
wire r5_297;
assign r5_297 = in[4]? r4_594 : r4_593;
wire r5_298;
assign r5_298 = in[4]? r4_596 : r4_595;
wire r5_299;
assign r5_299 = in[4]? r4_598 : r4_597;
wire r5_300;
assign r5_300 = in[4]? r4_600 : r4_599;
wire r5_301;
assign r5_301 = in[4]? r4_602 : r4_601;
wire r5_302;
assign r5_302 = in[4]? r4_604 : r4_603;
wire r5_303;
assign r5_303 = in[4]? r4_606 : r4_605;
wire r5_304;
assign r5_304 = in[4]? r4_608 : r4_607;
wire r5_305;
assign r5_305 = in[4]? r4_610 : r4_609;
wire r5_306;
assign r5_306 = in[4]? r4_612 : r4_611;
wire r5_307;
assign r5_307 = in[4]? r4_614 : r4_613;
wire r5_308;
assign r5_308 = in[4]? r4_616 : r4_615;
wire r5_309;
assign r5_309 = in[4]? r4_618 : r4_617;
wire r5_310;
assign r5_310 = in[4]? r4_620 : r4_619;
wire r5_311;
assign r5_311 = in[4]? r4_622 : r4_621;
wire r5_312;
assign r5_312 = in[4]? r4_624 : r4_623;
wire r5_313;
assign r5_313 = in[4]? r4_626 : r4_625;
wire r5_314;
assign r5_314 = in[4]? r4_628 : r4_627;
wire r5_315;
assign r5_315 = in[4]? r4_630 : r4_629;
wire r5_316;
assign r5_316 = in[4]? r4_632 : r4_631;
wire r5_317;
assign r5_317 = in[4]? r4_634 : r4_633;
wire r5_318;
assign r5_318 = in[4]? r4_636 : r4_635;
wire r5_319;
assign r5_319 = in[4]? r4_638 : r4_637;
wire r5_320;
assign r5_320 = in[4]? r4_640 : r4_639;
wire r5_321;
assign r5_321 = in[4]? r4_642 : r4_641;
wire r5_322;
assign r5_322 = in[4]? r4_644 : r4_643;
wire r5_323;
assign r5_323 = in[4]? r4_646 : r4_645;
wire r5_324;
assign r5_324 = in[4]? r4_648 : r4_647;
wire r5_325;
assign r5_325 = in[4]? r4_650 : r4_649;
wire r5_326;
assign r5_326 = in[4]? r4_652 : r4_651;
wire r5_327;
assign r5_327 = in[4]? r4_654 : r4_653;
wire r5_328;
assign r5_328 = in[4]? r4_656 : r4_655;
wire r5_329;
assign r5_329 = in[4]? r4_658 : r4_657;
wire r5_330;
assign r5_330 = in[4]? r4_660 : r4_659;
wire r5_331;
assign r5_331 = in[4]? r4_662 : r4_661;
wire r5_332;
assign r5_332 = in[4]? r4_664 : r4_663;
wire r5_333;
assign r5_333 = in[4]? r4_666 : r4_665;
wire r5_334;
assign r5_334 = in[4]? r4_668 : r4_667;
wire r5_335;
assign r5_335 = in[4]? r4_670 : r4_669;
wire r5_336;
assign r5_336 = in[4]? r4_672 : r4_671;
wire r5_337;
assign r5_337 = in[4]? r4_674 : r4_673;
wire r5_338;
assign r5_338 = in[4]? r4_676 : r4_675;
wire r5_339;
assign r5_339 = in[4]? r4_678 : r4_677;
wire r5_340;
assign r5_340 = in[4]? r4_680 : r4_679;
wire r5_341;
assign r5_341 = in[4]? r4_682 : r4_681;
wire r5_342;
assign r5_342 = in[4]? r4_684 : r4_683;
wire r5_343;
assign r5_343 = in[4]? r4_686 : r4_685;
wire r5_344;
assign r5_344 = in[4]? r4_688 : r4_687;
wire r5_345;
assign r5_345 = in[4]? r4_690 : r4_689;
wire r5_346;
assign r5_346 = in[4]? r4_692 : r4_691;
wire r5_347;
assign r5_347 = in[4]? r4_694 : r4_693;
wire r5_348;
assign r5_348 = in[4]? r4_696 : r4_695;
wire r5_349;
assign r5_349 = in[4]? r4_698 : r4_697;
wire r5_350;
assign r5_350 = in[4]? r4_700 : r4_699;
wire r5_351;
assign r5_351 = in[4]? r4_702 : r4_701;
wire r5_352;
assign r5_352 = in[4]? r4_704 : r4_703;
wire r5_353;
assign r5_353 = in[4]? r4_706 : r4_705;
wire r5_354;
assign r5_354 = in[4]? r4_708 : r4_707;
wire r5_355;
assign r5_355 = in[4]? r4_710 : r4_709;
wire r5_356;
assign r5_356 = in[4]? r4_712 : r4_711;
wire r5_357;
assign r5_357 = in[4]? r4_714 : r4_713;
wire r5_358;
assign r5_358 = in[4]? r4_716 : r4_715;
wire r5_359;
assign r5_359 = in[4]? r4_718 : r4_717;
wire r5_360;
assign r5_360 = in[4]? r4_720 : r4_719;
wire r5_361;
assign r5_361 = in[4]? r4_722 : r4_721;
wire r5_362;
assign r5_362 = in[4]? r4_724 : r4_723;
wire r5_363;
assign r5_363 = in[4]? r4_726 : r4_725;
wire r5_364;
assign r5_364 = in[4]? r4_728 : r4_727;
wire r5_365;
assign r5_365 = in[4]? r4_730 : r4_729;
wire r5_366;
assign r5_366 = in[4]? r4_732 : r4_731;
wire r5_367;
assign r5_367 = in[4]? r4_734 : r4_733;
wire r5_368;
assign r5_368 = in[4]? r4_736 : r4_735;
wire r5_369;
assign r5_369 = in[4]? r4_738 : r4_737;
wire r5_370;
assign r5_370 = in[4]? r4_740 : r4_739;
wire r5_371;
assign r5_371 = in[4]? r4_742 : r4_741;
wire r5_372;
assign r5_372 = in[4]? r4_744 : r4_743;
wire r5_373;
assign r5_373 = in[4]? r4_746 : r4_745;
wire r5_374;
assign r5_374 = in[4]? r4_748 : r4_747;
wire r5_375;
assign r5_375 = in[4]? r4_750 : r4_749;
wire r5_376;
assign r5_376 = in[4]? r4_752 : r4_751;
wire r5_377;
assign r5_377 = in[4]? r4_754 : r4_753;
wire r5_378;
assign r5_378 = in[4]? r4_756 : r4_755;
wire r5_379;
assign r5_379 = in[4]? r4_758 : r4_757;
wire r5_380;
assign r5_380 = in[4]? r4_760 : r4_759;
wire r5_381;
assign r5_381 = in[4]? r4_762 : r4_761;
wire r5_382;
assign r5_382 = in[4]? r4_764 : r4_763;
wire r5_383;
assign r5_383 = in[4]? r4_766 : r4_765;
wire r5_384;
assign r5_384 = in[4]? r4_768 : r4_767;
wire r5_385;
assign r5_385 = in[4]? r4_770 : r4_769;
wire r5_386;
assign r5_386 = in[4]? r4_772 : r4_771;
wire r5_387;
assign r5_387 = in[4]? r4_774 : r4_773;
wire r5_388;
assign r5_388 = in[4]? r4_776 : r4_775;
wire r5_389;
assign r5_389 = in[4]? r4_778 : r4_777;
wire r5_390;
assign r5_390 = in[4]? r4_780 : r4_779;
wire r5_391;
assign r5_391 = in[4]? r4_782 : r4_781;
wire r5_392;
assign r5_392 = in[4]? r4_784 : r4_783;
wire r5_393;
assign r5_393 = in[4]? r4_786 : r4_785;
wire r5_394;
assign r5_394 = in[4]? r4_788 : r4_787;
wire r5_395;
assign r5_395 = in[4]? r4_790 : r4_789;
wire r5_396;
assign r5_396 = in[4]? r4_792 : r4_791;
wire r5_397;
assign r5_397 = in[4]? r4_794 : r4_793;
wire r5_398;
assign r5_398 = in[4]? r4_796 : r4_795;
wire r5_399;
assign r5_399 = in[4]? r4_798 : r4_797;
wire r5_400;
assign r5_400 = in[4]? r4_800 : r4_799;
wire r5_401;
assign r5_401 = in[4]? r4_802 : r4_801;
wire r5_402;
assign r5_402 = in[4]? r4_804 : r4_803;
wire r5_403;
assign r5_403 = in[4]? r4_806 : r4_805;
wire r5_404;
assign r5_404 = in[4]? r4_808 : r4_807;
wire r5_405;
assign r5_405 = in[4]? r4_810 : r4_809;
wire r5_406;
assign r5_406 = in[4]? r4_812 : r4_811;
wire r5_407;
assign r5_407 = in[4]? r4_814 : r4_813;
wire r5_408;
assign r5_408 = in[4]? r4_816 : r4_815;
wire r5_409;
assign r5_409 = in[4]? r4_818 : r4_817;
wire r5_410;
assign r5_410 = in[4]? r4_820 : r4_819;
wire r5_411;
assign r5_411 = in[4]? r4_822 : r4_821;
wire r5_412;
assign r5_412 = in[4]? r4_824 : r4_823;
wire r5_413;
assign r5_413 = in[4]? r4_826 : r4_825;
wire r5_414;
assign r5_414 = in[4]? r4_828 : r4_827;
wire r5_415;
assign r5_415 = in[4]? r4_830 : r4_829;
wire r5_416;
assign r5_416 = in[4]? r4_832 : r4_831;
wire r5_417;
assign r5_417 = in[4]? r4_834 : r4_833;
wire r5_418;
assign r5_418 = in[4]? r4_836 : r4_835;
wire r5_419;
assign r5_419 = in[4]? r4_838 : r4_837;
wire r5_420;
assign r5_420 = in[4]? r4_840 : r4_839;
wire r5_421;
assign r5_421 = in[4]? r4_842 : r4_841;
wire r5_422;
assign r5_422 = in[4]? r4_844 : r4_843;
wire r5_423;
assign r5_423 = in[4]? r4_846 : r4_845;
wire r5_424;
assign r5_424 = in[4]? r4_848 : r4_847;
wire r5_425;
assign r5_425 = in[4]? r4_850 : r4_849;
wire r5_426;
assign r5_426 = in[4]? r4_852 : r4_851;
wire r5_427;
assign r5_427 = in[4]? r4_854 : r4_853;
wire r5_428;
assign r5_428 = in[4]? r4_856 : r4_855;
wire r5_429;
assign r5_429 = in[4]? r4_858 : r4_857;
wire r5_430;
assign r5_430 = in[4]? r4_860 : r4_859;
wire r5_431;
assign r5_431 = in[4]? r4_862 : r4_861;
wire r5_432;
assign r5_432 = in[4]? r4_864 : r4_863;
wire r5_433;
assign r5_433 = in[4]? r4_866 : r4_865;
wire r5_434;
assign r5_434 = in[4]? r4_868 : r4_867;
wire r5_435;
assign r5_435 = in[4]? r4_870 : r4_869;
wire r5_436;
assign r5_436 = in[4]? r4_872 : r4_871;
wire r5_437;
assign r5_437 = in[4]? r4_874 : r4_873;
wire r5_438;
assign r5_438 = in[4]? r4_876 : r4_875;
wire r5_439;
assign r5_439 = in[4]? r4_878 : r4_877;
wire r5_440;
assign r5_440 = in[4]? r4_880 : r4_879;
wire r5_441;
assign r5_441 = in[4]? r4_882 : r4_881;
wire r5_442;
assign r5_442 = in[4]? r4_884 : r4_883;
wire r5_443;
assign r5_443 = in[4]? r4_886 : r4_885;
wire r5_444;
assign r5_444 = in[4]? r4_888 : r4_887;
wire r5_445;
assign r5_445 = in[4]? r4_890 : r4_889;
wire r5_446;
assign r5_446 = in[4]? r4_892 : r4_891;
wire r5_447;
assign r5_447 = in[4]? r4_894 : r4_893;
wire r5_448;
assign r5_448 = in[4]? r4_896 : r4_895;
wire r5_449;
assign r5_449 = in[4]? r4_898 : r4_897;
wire r5_450;
assign r5_450 = in[4]? r4_900 : r4_899;
wire r5_451;
assign r5_451 = in[4]? r4_902 : r4_901;
wire r5_452;
assign r5_452 = in[4]? r4_904 : r4_903;
wire r5_453;
assign r5_453 = in[4]? r4_906 : r4_905;
wire r5_454;
assign r5_454 = in[4]? r4_908 : r4_907;
wire r5_455;
assign r5_455 = in[4]? r4_910 : r4_909;
wire r5_456;
assign r5_456 = in[4]? r4_912 : r4_911;
wire r5_457;
assign r5_457 = in[4]? r4_914 : r4_913;
wire r5_458;
assign r5_458 = in[4]? r4_916 : r4_915;
wire r5_459;
assign r5_459 = in[4]? r4_918 : r4_917;
wire r5_460;
assign r5_460 = in[4]? r4_920 : r4_919;
wire r5_461;
assign r5_461 = in[4]? r4_922 : r4_921;
wire r5_462;
assign r5_462 = in[4]? r4_924 : r4_923;
wire r5_463;
assign r5_463 = in[4]? r4_926 : r4_925;
wire r5_464;
assign r5_464 = in[4]? r4_928 : r4_927;
wire r5_465;
assign r5_465 = in[4]? r4_930 : r4_929;
wire r5_466;
assign r5_466 = in[4]? r4_932 : r4_931;
wire r5_467;
assign r5_467 = in[4]? r4_934 : r4_933;
wire r5_468;
assign r5_468 = in[4]? r4_936 : r4_935;
wire r5_469;
assign r5_469 = in[4]? r4_938 : r4_937;
wire r5_470;
assign r5_470 = in[4]? r4_940 : r4_939;
wire r5_471;
assign r5_471 = in[4]? r4_942 : r4_941;
wire r5_472;
assign r5_472 = in[4]? r4_944 : r4_943;
wire r5_473;
assign r5_473 = in[4]? r4_946 : r4_945;
wire r5_474;
assign r5_474 = in[4]? r4_948 : r4_947;
wire r5_475;
assign r5_475 = in[4]? r4_950 : r4_949;
wire r5_476;
assign r5_476 = in[4]? r4_952 : r4_951;
wire r5_477;
assign r5_477 = in[4]? r4_954 : r4_953;
wire r5_478;
assign r5_478 = in[4]? r4_956 : r4_955;
wire r5_479;
assign r5_479 = in[4]? r4_958 : r4_957;
wire r5_480;
assign r5_480 = in[4]? r4_960 : r4_959;
wire r5_481;
assign r5_481 = in[4]? r4_962 : r4_961;
wire r5_482;
assign r5_482 = in[4]? r4_964 : r4_963;
wire r5_483;
assign r5_483 = in[4]? r4_966 : r4_965;
wire r5_484;
assign r5_484 = in[4]? r4_968 : r4_967;
wire r5_485;
assign r5_485 = in[4]? r4_970 : r4_969;
wire r5_486;
assign r5_486 = in[4]? r4_972 : r4_971;
wire r5_487;
assign r5_487 = in[4]? r4_974 : r4_973;
wire r5_488;
assign r5_488 = in[4]? r4_976 : r4_975;
wire r5_489;
assign r5_489 = in[4]? r4_978 : r4_977;
wire r5_490;
assign r5_490 = in[4]? r4_980 : r4_979;
wire r5_491;
assign r5_491 = in[4]? r4_982 : r4_981;
wire r5_492;
assign r5_492 = in[4]? r4_984 : r4_983;
wire r5_493;
assign r5_493 = in[4]? r4_986 : r4_985;
wire r5_494;
assign r5_494 = in[4]? r4_988 : r4_987;
wire r5_495;
assign r5_495 = in[4]? r4_990 : r4_989;
wire r5_496;
assign r5_496 = in[4]? r4_992 : r4_991;
wire r5_497;
assign r5_497 = in[4]? r4_994 : r4_993;
wire r5_498;
assign r5_498 = in[4]? r4_996 : r4_995;
wire r5_499;
assign r5_499 = in[4]? r4_998 : r4_997;
wire r5_500;
assign r5_500 = in[4]? r4_1000 : r4_999;
wire r5_501;
assign r5_501 = in[4]? r4_1002 : r4_1001;
wire r5_502;
assign r5_502 = in[4]? r4_1004 : r4_1003;
wire r5_503;
assign r5_503 = in[4]? r4_1006 : r4_1005;
wire r5_504;
assign r5_504 = in[4]? r4_1008 : r4_1007;
wire r5_505;
assign r5_505 = in[4]? r4_1010 : r4_1009;
wire r5_506;
assign r5_506 = in[4]? r4_1012 : r4_1011;
wire r5_507;
assign r5_507 = in[4]? r4_1014 : r4_1013;
wire r5_508;
assign r5_508 = in[4]? r4_1016 : r4_1015;
wire r5_509;
assign r5_509 = in[4]? r4_1018 : r4_1017;
wire r5_510;
assign r5_510 = in[4]? r4_1020 : r4_1019;
wire r5_511;
assign r5_511 = in[4]? r4_1022 : r4_1021;
wire r5_512;
assign r5_512 = in[4]? r4_1024 : r4_1023;
wire r5_513;
assign r5_513 = in[4]? r4_1026 : r4_1025;
wire r5_514;
assign r5_514 = in[4]? r4_1028 : r4_1027;
wire r5_515;
assign r5_515 = in[4]? r4_1030 : r4_1029;
wire r5_516;
assign r5_516 = in[4]? r4_1032 : r4_1031;
wire r5_517;
assign r5_517 = in[4]? r4_1034 : r4_1033;
wire r5_518;
assign r5_518 = in[4]? r4_1036 : r4_1035;
wire r5_519;
assign r5_519 = in[4]? r4_1038 : r4_1037;
wire r5_520;
assign r5_520 = in[4]? r4_1040 : r4_1039;
wire r5_521;
assign r5_521 = in[4]? r4_1042 : r4_1041;
wire r5_522;
assign r5_522 = in[4]? r4_1044 : r4_1043;
wire r5_523;
assign r5_523 = in[4]? r4_1046 : r4_1045;
wire r5_524;
assign r5_524 = in[4]? r4_1048 : r4_1047;
wire r5_525;
assign r5_525 = in[4]? r4_1050 : r4_1049;
wire r5_526;
assign r5_526 = in[4]? r4_1052 : r4_1051;
wire r5_527;
assign r5_527 = in[4]? r4_1054 : r4_1053;
wire r5_528;
assign r5_528 = in[4]? r4_1056 : r4_1055;
wire r5_529;
assign r5_529 = in[4]? r4_1058 : r4_1057;
wire r5_530;
assign r5_530 = in[4]? r4_1060 : r4_1059;
wire r5_531;
assign r5_531 = in[4]? r4_1062 : r4_1061;
wire r5_532;
assign r5_532 = in[4]? r4_1064 : r4_1063;
wire r5_533;
assign r5_533 = in[4]? r4_1066 : r4_1065;
wire r5_534;
assign r5_534 = in[4]? r4_1068 : r4_1067;
wire r5_535;
assign r5_535 = in[4]? r4_1070 : r4_1069;
wire r5_536;
assign r5_536 = in[4]? r4_1072 : r4_1071;
wire r5_537;
assign r5_537 = in[4]? r4_1074 : r4_1073;
wire r5_538;
assign r5_538 = in[4]? r4_1076 : r4_1075;
wire r5_539;
assign r5_539 = in[4]? r4_1078 : r4_1077;
wire r5_540;
assign r5_540 = in[4]? r4_1080 : r4_1079;
wire r5_541;
assign r5_541 = in[4]? r4_1082 : r4_1081;
wire r5_542;
assign r5_542 = in[4]? r4_1084 : r4_1083;
wire r5_543;
assign r5_543 = in[4]? r4_1086 : r4_1085;
wire r5_544;
assign r5_544 = in[4]? r4_1088 : r4_1087;
wire r5_545;
assign r5_545 = in[4]? r4_1090 : r4_1089;
wire r5_546;
assign r5_546 = in[4]? r4_1092 : r4_1091;
wire r5_547;
assign r5_547 = in[4]? r4_1094 : r4_1093;
wire r5_548;
assign r5_548 = in[4]? r4_1096 : r4_1095;
wire r5_549;
assign r5_549 = in[4]? r4_1098 : r4_1097;
wire r5_550;
assign r5_550 = in[4]? r4_1100 : r4_1099;
wire r5_551;
assign r5_551 = in[4]? r4_1102 : r4_1101;
wire r5_552;
assign r5_552 = in[4]? r4_1104 : r4_1103;
wire r5_553;
assign r5_553 = in[4]? r4_1106 : r4_1105;
wire r5_554;
assign r5_554 = in[4]? r4_1108 : r4_1107;
wire r5_555;
assign r5_555 = in[4]? r4_1110 : r4_1109;
wire r5_556;
assign r5_556 = in[4]? r4_1112 : r4_1111;
wire r5_557;
assign r5_557 = in[4]? r4_1114 : r4_1113;
wire r5_558;
assign r5_558 = in[4]? r4_1116 : r4_1115;
wire r5_559;
assign r5_559 = in[4]? r4_1118 : r4_1117;
wire r5_560;
assign r5_560 = in[4]? r4_1120 : r4_1119;
wire r5_561;
assign r5_561 = in[4]? r4_1122 : r4_1121;
wire r5_562;
assign r5_562 = in[4]? r4_1124 : r4_1123;
wire r5_563;
assign r5_563 = in[4]? r4_1126 : r4_1125;
wire r5_564;
assign r5_564 = in[4]? r4_1128 : r4_1127;
wire r5_565;
assign r5_565 = in[4]? r4_1130 : r4_1129;
wire r5_566;
assign r5_566 = in[4]? r4_1132 : r4_1131;
wire r5_567;
assign r5_567 = in[4]? r4_1134 : r4_1133;
wire r5_568;
assign r5_568 = in[4]? r4_1136 : r4_1135;
wire r5_569;
assign r5_569 = in[4]? r4_1138 : r4_1137;
wire r5_570;
assign r5_570 = in[4]? r4_1140 : r4_1139;
wire r5_571;
assign r5_571 = in[4]? r4_1142 : r4_1141;
wire r5_572;
assign r5_572 = in[4]? r4_1144 : r4_1143;
wire r5_573;
assign r5_573 = in[4]? r4_1146 : r4_1145;
wire r5_574;
assign r5_574 = in[4]? r4_1148 : r4_1147;
wire r5_575;
assign r5_575 = in[4]? r4_1150 : r4_1149;
wire r5_576;
assign r5_576 = in[4]? r4_1152 : r4_1151;
wire r5_577;
assign r5_577 = in[4]? r4_1154 : r4_1153;
wire r5_578;
assign r5_578 = in[4]? r4_1156 : r4_1155;
wire r5_579;
assign r5_579 = in[4]? r4_1158 : r4_1157;
wire r5_580;
assign r5_580 = in[4]? r4_1160 : r4_1159;
wire r5_581;
assign r5_581 = in[4]? r4_1162 : r4_1161;
wire r5_582;
assign r5_582 = in[4]? r4_1164 : r4_1163;
wire r5_583;
assign r5_583 = in[4]? r4_1166 : r4_1165;
wire r5_584;
assign r5_584 = in[4]? r4_1168 : r4_1167;
wire r5_585;
assign r5_585 = in[4]? r4_1170 : r4_1169;
wire r5_586;
assign r5_586 = in[4]? r4_1172 : r4_1171;
wire r5_587;
assign r5_587 = in[4]? r4_1174 : r4_1173;
wire r5_588;
assign r5_588 = in[4]? r4_1176 : r4_1175;
wire r5_589;
assign r5_589 = in[4]? r4_1178 : r4_1177;
wire r5_590;
assign r5_590 = in[4]? r4_1180 : r4_1179;
wire r5_591;
assign r5_591 = in[4]? r4_1182 : r4_1181;
wire r5_592;
assign r5_592 = in[4]? r4_1184 : r4_1183;
wire r5_593;
assign r5_593 = in[4]? r4_1186 : r4_1185;
wire r5_594;
assign r5_594 = in[4]? r4_1188 : r4_1187;
wire r5_595;
assign r5_595 = in[4]? r4_1190 : r4_1189;
wire r5_596;
assign r5_596 = in[4]? r4_1192 : r4_1191;
wire r5_597;
assign r5_597 = in[4]? r4_1194 : r4_1193;
wire r5_598;
assign r5_598 = in[4]? r4_1196 : r4_1195;
wire r5_599;
assign r5_599 = in[4]? r4_1198 : r4_1197;
wire r5_600;
assign r5_600 = in[4]? r4_1200 : r4_1199;
wire r5_601;
assign r5_601 = in[4]? r4_1202 : r4_1201;
wire r5_602;
assign r5_602 = in[4]? r4_1204 : r4_1203;
wire r5_603;
assign r5_603 = in[4]? r4_1206 : r4_1205;
wire r5_604;
assign r5_604 = in[4]? r4_1208 : r4_1207;
wire r5_605;
assign r5_605 = in[4]? r4_1210 : r4_1209;
wire r5_606;
assign r5_606 = in[4]? r4_1212 : r4_1211;
wire r5_607;
assign r5_607 = in[4]? r4_1214 : r4_1213;
wire r5_608;
assign r5_608 = in[4]? r4_1216 : r4_1215;
wire r5_609;
assign r5_609 = in[4]? r4_1218 : r4_1217;
wire r5_610;
assign r5_610 = in[4]? r4_1220 : r4_1219;
wire r5_611;
assign r5_611 = in[4]? r4_1222 : r4_1221;
wire r5_612;
assign r5_612 = in[4]? r4_1224 : r4_1223;
wire r5_613;
assign r5_613 = in[4]? r4_1226 : r4_1225;
wire r5_614;
assign r5_614 = in[4]? r4_1228 : r4_1227;
wire r5_615;
assign r5_615 = in[4]? r4_1230 : r4_1229;
wire r5_616;
assign r5_616 = in[4]? r4_1232 : r4_1231;
wire r5_617;
assign r5_617 = in[4]? r4_1234 : r4_1233;
wire r5_618;
assign r5_618 = in[4]? r4_1236 : r4_1235;
wire r5_619;
assign r5_619 = in[4]? r4_1238 : r4_1237;
wire r5_620;
assign r5_620 = in[4]? r4_1240 : r4_1239;
wire r5_621;
assign r5_621 = in[4]? r4_1242 : r4_1241;
wire r5_622;
assign r5_622 = in[4]? r4_1244 : r4_1243;
wire r5_623;
assign r5_623 = in[4]? r4_1246 : r4_1245;
wire r5_624;
assign r5_624 = in[4]? r4_1248 : r4_1247;
wire r5_625;
assign r5_625 = in[4]? r4_1250 : r4_1249;
wire r5_626;
assign r5_626 = in[4]? r4_1252 : r4_1251;
wire r5_627;
assign r5_627 = in[4]? r4_1254 : r4_1253;
wire r5_628;
assign r5_628 = in[4]? r4_1256 : r4_1255;
wire r5_629;
assign r5_629 = in[4]? r4_1258 : r4_1257;
wire r5_630;
assign r5_630 = in[4]? r4_1260 : r4_1259;
wire r5_631;
assign r5_631 = in[4]? r4_1262 : r4_1261;
wire r5_632;
assign r5_632 = in[4]? r4_1264 : r4_1263;
wire r5_633;
assign r5_633 = in[4]? r4_1266 : r4_1265;
wire r5_634;
assign r5_634 = in[4]? r4_1268 : r4_1267;
wire r5_635;
assign r5_635 = in[4]? r4_1270 : r4_1269;
wire r5_636;
assign r5_636 = in[4]? r4_1272 : r4_1271;
wire r5_637;
assign r5_637 = in[4]? r4_1274 : r4_1273;
wire r5_638;
assign r5_638 = in[4]? r4_1276 : r4_1275;
wire r5_639;
assign r5_639 = in[4]? r4_1278 : r4_1277;
wire r5_640;
assign r5_640 = in[4]? r4_1280 : r4_1279;
wire r5_641;
assign r5_641 = in[4]? r4_1282 : r4_1281;
wire r5_642;
assign r5_642 = in[4]? r4_1284 : r4_1283;
wire r6_1;
assign r6_1 = in[5]? r5_2 : r5_1;
wire r6_2;
assign r6_2 = in[5]? r5_4 : r5_3;
wire r6_3;
assign r6_3 = in[5]? r5_6 : r5_5;
wire r6_4;
assign r6_4 = in[5]? r5_8 : r5_7;
wire r6_5;
assign r6_5 = in[5]? r5_10 : r5_9;
wire r6_6;
assign r6_6 = in[5]? r5_12 : r5_11;
wire r6_7;
assign r6_7 = in[5]? r5_14 : r5_13;
wire r6_8;
assign r6_8 = in[5]? r5_16 : r5_15;
wire r6_9;
assign r6_9 = in[5]? r5_18 : r5_17;
wire r6_10;
assign r6_10 = in[5]? r5_20 : r5_19;
wire r6_11;
assign r6_11 = in[5]? r5_22 : r5_21;
wire r6_12;
assign r6_12 = in[5]? r5_24 : r5_23;
wire r6_13;
assign r6_13 = in[5]? r5_26 : r5_25;
wire r6_14;
assign r6_14 = in[5]? r5_28 : r5_27;
wire r6_15;
assign r6_15 = in[5]? r5_30 : r5_29;
wire r6_16;
assign r6_16 = in[5]? r5_32 : r5_31;
wire r6_17;
assign r6_17 = in[5]? r5_34 : r5_33;
wire r6_18;
assign r6_18 = in[5]? r5_36 : r5_35;
wire r6_19;
assign r6_19 = in[5]? r5_38 : r5_37;
wire r6_20;
assign r6_20 = in[5]? r5_40 : r5_39;
wire r6_21;
assign r6_21 = in[5]? r5_42 : r5_41;
wire r6_22;
assign r6_22 = in[5]? r5_44 : r5_43;
wire r6_23;
assign r6_23 = in[5]? r5_46 : r5_45;
wire r6_24;
assign r6_24 = in[5]? r5_48 : r5_47;
wire r6_25;
assign r6_25 = in[5]? r5_50 : r5_49;
wire r6_26;
assign r6_26 = in[5]? r5_52 : r5_51;
wire r6_27;
assign r6_27 = in[5]? r5_54 : r5_53;
wire r6_28;
assign r6_28 = in[5]? r5_56 : r5_55;
wire r6_29;
assign r6_29 = in[5]? r5_58 : r5_57;
wire r6_30;
assign r6_30 = in[5]? r5_60 : r5_59;
wire r6_31;
assign r6_31 = in[5]? r5_62 : r5_61;
wire r6_32;
assign r6_32 = in[5]? r5_64 : r5_63;
wire r6_33;
assign r6_33 = in[5]? r5_66 : r5_65;
wire r6_34;
assign r6_34 = in[5]? r5_68 : r5_67;
wire r6_35;
assign r6_35 = in[5]? r5_70 : r5_69;
wire r6_36;
assign r6_36 = in[5]? r5_72 : r5_71;
wire r6_37;
assign r6_37 = in[5]? r5_74 : r5_73;
wire r6_38;
assign r6_38 = in[5]? r5_76 : r5_75;
wire r6_39;
assign r6_39 = in[5]? r5_78 : r5_77;
wire r6_40;
assign r6_40 = in[5]? r5_80 : r5_79;
wire r6_41;
assign r6_41 = in[5]? r5_82 : r5_81;
wire r6_42;
assign r6_42 = in[5]? r5_84 : r5_83;
wire r6_43;
assign r6_43 = in[5]? r5_86 : r5_85;
wire r6_44;
assign r6_44 = in[5]? r5_88 : r5_87;
wire r6_45;
assign r6_45 = in[5]? r5_90 : r5_89;
wire r6_46;
assign r6_46 = in[5]? r5_92 : r5_91;
wire r6_47;
assign r6_47 = in[5]? r5_94 : r5_93;
wire r6_48;
assign r6_48 = in[5]? r5_96 : r5_95;
wire r6_49;
assign r6_49 = in[5]? r5_98 : r5_97;
wire r6_50;
assign r6_50 = in[5]? r5_100 : r5_99;
wire r6_51;
assign r6_51 = in[5]? r5_102 : r5_101;
wire r6_52;
assign r6_52 = in[5]? r5_104 : r5_103;
wire r6_53;
assign r6_53 = in[5]? r5_106 : r5_105;
wire r6_54;
assign r6_54 = in[5]? r5_108 : r5_107;
wire r6_55;
assign r6_55 = in[5]? r5_110 : r5_109;
wire r6_56;
assign r6_56 = in[5]? r5_112 : r5_111;
wire r6_57;
assign r6_57 = in[5]? r5_114 : r5_113;
wire r6_58;
assign r6_58 = in[5]? r5_116 : r5_115;
wire r6_59;
assign r6_59 = in[5]? r5_118 : r5_117;
wire r6_60;
assign r6_60 = in[5]? r5_120 : r5_119;
wire r6_61;
assign r6_61 = in[5]? r5_122 : r5_121;
wire r6_62;
assign r6_62 = in[5]? r5_124 : r5_123;
wire r6_63;
assign r6_63 = in[5]? r5_126 : r5_125;
wire r6_64;
assign r6_64 = in[5]? r5_128 : r5_127;
wire r6_65;
assign r6_65 = in[5]? r5_130 : r5_129;
wire r6_66;
assign r6_66 = in[5]? r5_132 : r5_131;
wire r6_67;
assign r6_67 = in[5]? r5_134 : r5_133;
wire r6_68;
assign r6_68 = in[5]? r5_136 : r5_135;
wire r6_69;
assign r6_69 = in[5]? r5_138 : r5_137;
wire r6_70;
assign r6_70 = in[5]? r5_140 : r5_139;
wire r6_71;
assign r6_71 = in[5]? r5_142 : r5_141;
wire r6_72;
assign r6_72 = in[5]? r5_144 : r5_143;
wire r6_73;
assign r6_73 = in[5]? r5_146 : r5_145;
wire r6_74;
assign r6_74 = in[5]? r5_148 : r5_147;
wire r6_75;
assign r6_75 = in[5]? r5_150 : r5_149;
wire r6_76;
assign r6_76 = in[5]? r5_152 : r5_151;
wire r6_77;
assign r6_77 = in[5]? r5_154 : r5_153;
wire r6_78;
assign r6_78 = in[5]? r5_156 : r5_155;
wire r6_79;
assign r6_79 = in[5]? r5_158 : r5_157;
wire r6_80;
assign r6_80 = in[5]? r5_160 : r5_159;
wire r6_81;
assign r6_81 = in[5]? r5_162 : r5_161;
wire r6_82;
assign r6_82 = in[5]? r5_164 : r5_163;
wire r6_83;
assign r6_83 = in[5]? r5_166 : r5_165;
wire r6_84;
assign r6_84 = in[5]? r5_168 : r5_167;
wire r6_85;
assign r6_85 = in[5]? r5_170 : r5_169;
wire r6_86;
assign r6_86 = in[5]? r5_172 : r5_171;
wire r6_87;
assign r6_87 = in[5]? r5_174 : r5_173;
wire r6_88;
assign r6_88 = in[5]? r5_176 : r5_175;
wire r6_89;
assign r6_89 = in[5]? r5_178 : r5_177;
wire r6_90;
assign r6_90 = in[5]? r5_180 : r5_179;
wire r6_91;
assign r6_91 = in[5]? r5_182 : r5_181;
wire r6_92;
assign r6_92 = in[5]? r5_184 : r5_183;
wire r6_93;
assign r6_93 = in[5]? r5_186 : r5_185;
wire r6_94;
assign r6_94 = in[5]? r5_188 : r5_187;
wire r6_95;
assign r6_95 = in[5]? r5_190 : r5_189;
wire r6_96;
assign r6_96 = in[5]? r5_192 : r5_191;
wire r6_97;
assign r6_97 = in[5]? r5_194 : r5_193;
wire r6_98;
assign r6_98 = in[5]? r5_196 : r5_195;
wire r6_99;
assign r6_99 = in[5]? r5_198 : r5_197;
wire r6_100;
assign r6_100 = in[5]? r5_200 : r5_199;
wire r6_101;
assign r6_101 = in[5]? r5_202 : r5_201;
wire r6_102;
assign r6_102 = in[5]? r5_204 : r5_203;
wire r6_103;
assign r6_103 = in[5]? r5_206 : r5_205;
wire r6_104;
assign r6_104 = in[5]? r5_208 : r5_207;
wire r6_105;
assign r6_105 = in[5]? r5_210 : r5_209;
wire r6_106;
assign r6_106 = in[5]? r5_212 : r5_211;
wire r6_107;
assign r6_107 = in[5]? r5_214 : r5_213;
wire r6_108;
assign r6_108 = in[5]? r5_216 : r5_215;
wire r6_109;
assign r6_109 = in[5]? r5_218 : r5_217;
wire r6_110;
assign r6_110 = in[5]? r5_220 : r5_219;
wire r6_111;
assign r6_111 = in[5]? r5_222 : r5_221;
wire r6_112;
assign r6_112 = in[5]? r5_224 : r5_223;
wire r6_113;
assign r6_113 = in[5]? r5_226 : r5_225;
wire r6_114;
assign r6_114 = in[5]? r5_228 : r5_227;
wire r6_115;
assign r6_115 = in[5]? r5_230 : r5_229;
wire r6_116;
assign r6_116 = in[5]? r5_232 : r5_231;
wire r6_117;
assign r6_117 = in[5]? r5_234 : r5_233;
wire r6_118;
assign r6_118 = in[5]? r5_236 : r5_235;
wire r6_119;
assign r6_119 = in[5]? r5_238 : r5_237;
wire r6_120;
assign r6_120 = in[5]? r5_240 : r5_239;
wire r6_121;
assign r6_121 = in[5]? r5_242 : r5_241;
wire r6_122;
assign r6_122 = in[5]? r5_244 : r5_243;
wire r6_123;
assign r6_123 = in[5]? r5_246 : r5_245;
wire r6_124;
assign r6_124 = in[5]? r5_248 : r5_247;
wire r6_125;
assign r6_125 = in[5]? r5_250 : r5_249;
wire r6_126;
assign r6_126 = in[5]? r5_252 : r5_251;
wire r6_127;
assign r6_127 = in[5]? r5_254 : r5_253;
wire r6_128;
assign r6_128 = in[5]? r5_256 : r5_255;
wire r6_129;
assign r6_129 = in[5]? r5_258 : r5_257;
wire r6_130;
assign r6_130 = in[5]? r5_260 : r5_259;
wire r6_131;
assign r6_131 = in[5]? r5_262 : r5_261;
wire r6_132;
assign r6_132 = in[5]? r5_264 : r5_263;
wire r6_133;
assign r6_133 = in[5]? r5_266 : r5_265;
wire r6_134;
assign r6_134 = in[5]? r5_268 : r5_267;
wire r6_135;
assign r6_135 = in[5]? r5_270 : r5_269;
wire r6_136;
assign r6_136 = in[5]? r5_272 : r5_271;
wire r6_137;
assign r6_137 = in[5]? r5_274 : r5_273;
wire r6_138;
assign r6_138 = in[5]? r5_276 : r5_275;
wire r6_139;
assign r6_139 = in[5]? r5_278 : r5_277;
wire r6_140;
assign r6_140 = in[5]? r5_280 : r5_279;
wire r6_141;
assign r6_141 = in[5]? r5_282 : r5_281;
wire r6_142;
assign r6_142 = in[5]? r5_284 : r5_283;
wire r6_143;
assign r6_143 = in[5]? r5_286 : r5_285;
wire r6_144;
assign r6_144 = in[5]? r5_288 : r5_287;
wire r6_145;
assign r6_145 = in[5]? r5_290 : r5_289;
wire r6_146;
assign r6_146 = in[5]? r5_292 : r5_291;
wire r6_147;
assign r6_147 = in[5]? r5_294 : r5_293;
wire r6_148;
assign r6_148 = in[5]? r5_296 : r5_295;
wire r6_149;
assign r6_149 = in[5]? r5_298 : r5_297;
wire r6_150;
assign r6_150 = in[5]? r5_300 : r5_299;
wire r6_151;
assign r6_151 = in[5]? r5_302 : r5_301;
wire r6_152;
assign r6_152 = in[5]? r5_304 : r5_303;
wire r6_153;
assign r6_153 = in[5]? r5_306 : r5_305;
wire r6_154;
assign r6_154 = in[5]? r5_308 : r5_307;
wire r6_155;
assign r6_155 = in[5]? r5_310 : r5_309;
wire r6_156;
assign r6_156 = in[5]? r5_312 : r5_311;
wire r6_157;
assign r6_157 = in[5]? r5_314 : r5_313;
wire r6_158;
assign r6_158 = in[5]? r5_316 : r5_315;
wire r6_159;
assign r6_159 = in[5]? r5_318 : r5_317;
wire r6_160;
assign r6_160 = in[5]? r5_320 : r5_319;
wire r6_161;
assign r6_161 = in[5]? r5_322 : r5_321;
wire r6_162;
assign r6_162 = in[5]? r5_324 : r5_323;
wire r6_163;
assign r6_163 = in[5]? r5_326 : r5_325;
wire r6_164;
assign r6_164 = in[5]? r5_328 : r5_327;
wire r6_165;
assign r6_165 = in[5]? r5_330 : r5_329;
wire r6_166;
assign r6_166 = in[5]? r5_332 : r5_331;
wire r6_167;
assign r6_167 = in[5]? r5_334 : r5_333;
wire r6_168;
assign r6_168 = in[5]? r5_336 : r5_335;
wire r6_169;
assign r6_169 = in[5]? r5_338 : r5_337;
wire r6_170;
assign r6_170 = in[5]? r5_340 : r5_339;
wire r6_171;
assign r6_171 = in[5]? r5_342 : r5_341;
wire r6_172;
assign r6_172 = in[5]? r5_344 : r5_343;
wire r6_173;
assign r6_173 = in[5]? r5_346 : r5_345;
wire r6_174;
assign r6_174 = in[5]? r5_348 : r5_347;
wire r6_175;
assign r6_175 = in[5]? r5_350 : r5_349;
wire r6_176;
assign r6_176 = in[5]? r5_352 : r5_351;
wire r6_177;
assign r6_177 = in[5]? r5_354 : r5_353;
wire r6_178;
assign r6_178 = in[5]? r5_356 : r5_355;
wire r6_179;
assign r6_179 = in[5]? r5_358 : r5_357;
wire r6_180;
assign r6_180 = in[5]? r5_360 : r5_359;
wire r6_181;
assign r6_181 = in[5]? r5_362 : r5_361;
wire r6_182;
assign r6_182 = in[5]? r5_364 : r5_363;
wire r6_183;
assign r6_183 = in[5]? r5_366 : r5_365;
wire r6_184;
assign r6_184 = in[5]? r5_368 : r5_367;
wire r6_185;
assign r6_185 = in[5]? r5_370 : r5_369;
wire r6_186;
assign r6_186 = in[5]? r5_372 : r5_371;
wire r6_187;
assign r6_187 = in[5]? r5_374 : r5_373;
wire r6_188;
assign r6_188 = in[5]? r5_376 : r5_375;
wire r6_189;
assign r6_189 = in[5]? r5_378 : r5_377;
wire r6_190;
assign r6_190 = in[5]? r5_380 : r5_379;
wire r6_191;
assign r6_191 = in[5]? r5_382 : r5_381;
wire r6_192;
assign r6_192 = in[5]? r5_384 : r5_383;
wire r6_193;
assign r6_193 = in[5]? r5_386 : r5_385;
wire r6_194;
assign r6_194 = in[5]? r5_388 : r5_387;
wire r6_195;
assign r6_195 = in[5]? r5_390 : r5_389;
wire r6_196;
assign r6_196 = in[5]? r5_392 : r5_391;
wire r6_197;
assign r6_197 = in[5]? r5_394 : r5_393;
wire r6_198;
assign r6_198 = in[5]? r5_396 : r5_395;
wire r6_199;
assign r6_199 = in[5]? r5_398 : r5_397;
wire r6_200;
assign r6_200 = in[5]? r5_400 : r5_399;
wire r6_201;
assign r6_201 = in[5]? r5_402 : r5_401;
wire r6_202;
assign r6_202 = in[5]? r5_404 : r5_403;
wire r6_203;
assign r6_203 = in[5]? r5_406 : r5_405;
wire r6_204;
assign r6_204 = in[5]? r5_408 : r5_407;
wire r6_205;
assign r6_205 = in[5]? r5_410 : r5_409;
wire r6_206;
assign r6_206 = in[5]? r5_412 : r5_411;
wire r6_207;
assign r6_207 = in[5]? r5_414 : r5_413;
wire r6_208;
assign r6_208 = in[5]? r5_416 : r5_415;
wire r6_209;
assign r6_209 = in[5]? r5_418 : r5_417;
wire r6_210;
assign r6_210 = in[5]? r5_420 : r5_419;
wire r6_211;
assign r6_211 = in[5]? r5_422 : r5_421;
wire r6_212;
assign r6_212 = in[5]? r5_424 : r5_423;
wire r6_213;
assign r6_213 = in[5]? r5_426 : r5_425;
wire r6_214;
assign r6_214 = in[5]? r5_428 : r5_427;
wire r6_215;
assign r6_215 = in[5]? r5_430 : r5_429;
wire r6_216;
assign r6_216 = in[5]? r5_432 : r5_431;
wire r6_217;
assign r6_217 = in[5]? r5_434 : r5_433;
wire r6_218;
assign r6_218 = in[5]? r5_436 : r5_435;
wire r6_219;
assign r6_219 = in[5]? r5_438 : r5_437;
wire r6_220;
assign r6_220 = in[5]? r5_440 : r5_439;
wire r6_221;
assign r6_221 = in[5]? r5_442 : r5_441;
wire r6_222;
assign r6_222 = in[5]? r5_444 : r5_443;
wire r6_223;
assign r6_223 = in[5]? r5_446 : r5_445;
wire r6_224;
assign r6_224 = in[5]? r5_448 : r5_447;
wire r6_225;
assign r6_225 = in[5]? r5_450 : r5_449;
wire r6_226;
assign r6_226 = in[5]? r5_452 : r5_451;
wire r6_227;
assign r6_227 = in[5]? r5_454 : r5_453;
wire r6_228;
assign r6_228 = in[5]? r5_456 : r5_455;
wire r6_229;
assign r6_229 = in[5]? r5_458 : r5_457;
wire r6_230;
assign r6_230 = in[5]? r5_460 : r5_459;
wire r6_231;
assign r6_231 = in[5]? r5_462 : r5_461;
wire r6_232;
assign r6_232 = in[5]? r5_464 : r5_463;
wire r6_233;
assign r6_233 = in[5]? r5_466 : r5_465;
wire r6_234;
assign r6_234 = in[5]? r5_468 : r5_467;
wire r6_235;
assign r6_235 = in[5]? r5_470 : r5_469;
wire r6_236;
assign r6_236 = in[5]? r5_472 : r5_471;
wire r6_237;
assign r6_237 = in[5]? r5_474 : r5_473;
wire r6_238;
assign r6_238 = in[5]? r5_476 : r5_475;
wire r6_239;
assign r6_239 = in[5]? r5_478 : r5_477;
wire r6_240;
assign r6_240 = in[5]? r5_480 : r5_479;
wire r6_241;
assign r6_241 = in[5]? r5_482 : r5_481;
wire r6_242;
assign r6_242 = in[5]? r5_484 : r5_483;
wire r6_243;
assign r6_243 = in[5]? r5_486 : r5_485;
wire r6_244;
assign r6_244 = in[5]? r5_488 : r5_487;
wire r6_245;
assign r6_245 = in[5]? r5_490 : r5_489;
wire r6_246;
assign r6_246 = in[5]? r5_492 : r5_491;
wire r6_247;
assign r6_247 = in[5]? r5_494 : r5_493;
wire r6_248;
assign r6_248 = in[5]? r5_496 : r5_495;
wire r6_249;
assign r6_249 = in[5]? r5_498 : r5_497;
wire r6_250;
assign r6_250 = in[5]? r5_500 : r5_499;
wire r6_251;
assign r6_251 = in[5]? r5_502 : r5_501;
wire r6_252;
assign r6_252 = in[5]? r5_504 : r5_503;
wire r6_253;
assign r6_253 = in[5]? r5_506 : r5_505;
wire r6_254;
assign r6_254 = in[5]? r5_508 : r5_507;
wire r6_255;
assign r6_255 = in[5]? r5_510 : r5_509;
wire r6_256;
assign r6_256 = in[5]? r5_512 : r5_511;
wire r6_257;
assign r6_257 = in[5]? r5_514 : r5_513;
wire r6_258;
assign r6_258 = in[5]? r5_516 : r5_515;
wire r6_259;
assign r6_259 = in[5]? r5_518 : r5_517;
wire r6_260;
assign r6_260 = in[5]? r5_520 : r5_519;
wire r6_261;
assign r6_261 = in[5]? r5_522 : r5_521;
wire r6_262;
assign r6_262 = in[5]? r5_524 : r5_523;
wire r6_263;
assign r6_263 = in[5]? r5_526 : r5_525;
wire r6_264;
assign r6_264 = in[5]? r5_528 : r5_527;
wire r6_265;
assign r6_265 = in[5]? r5_530 : r5_529;
wire r6_266;
assign r6_266 = in[5]? r5_532 : r5_531;
wire r6_267;
assign r6_267 = in[5]? r5_534 : r5_533;
wire r6_268;
assign r6_268 = in[5]? r5_536 : r5_535;
wire r6_269;
assign r6_269 = in[5]? r5_538 : r5_537;
wire r6_270;
assign r6_270 = in[5]? r5_540 : r5_539;
wire r6_271;
assign r6_271 = in[5]? r5_542 : r5_541;
wire r6_272;
assign r6_272 = in[5]? r5_544 : r5_543;
wire r6_273;
assign r6_273 = in[5]? r5_546 : r5_545;
wire r6_274;
assign r6_274 = in[5]? r5_548 : r5_547;
wire r6_275;
assign r6_275 = in[5]? r5_550 : r5_549;
wire r6_276;
assign r6_276 = in[5]? r5_552 : r5_551;
wire r6_277;
assign r6_277 = in[5]? r5_554 : r5_553;
wire r6_278;
assign r6_278 = in[5]? r5_556 : r5_555;
wire r6_279;
assign r6_279 = in[5]? r5_558 : r5_557;
wire r6_280;
assign r6_280 = in[5]? r5_560 : r5_559;
wire r6_281;
assign r6_281 = in[5]? r5_562 : r5_561;
wire r6_282;
assign r6_282 = in[5]? r5_564 : r5_563;
wire r6_283;
assign r6_283 = in[5]? r5_566 : r5_565;
wire r6_284;
assign r6_284 = in[5]? r5_568 : r5_567;
wire r6_285;
assign r6_285 = in[5]? r5_570 : r5_569;
wire r6_286;
assign r6_286 = in[5]? r5_572 : r5_571;
wire r6_287;
assign r6_287 = in[5]? r5_574 : r5_573;
wire r6_288;
assign r6_288 = in[5]? r5_576 : r5_575;
wire r6_289;
assign r6_289 = in[5]? r5_578 : r5_577;
wire r6_290;
assign r6_290 = in[5]? r5_580 : r5_579;
wire r6_291;
assign r6_291 = in[5]? r5_582 : r5_581;
wire r6_292;
assign r6_292 = in[5]? r5_584 : r5_583;
wire r6_293;
assign r6_293 = in[5]? r5_586 : r5_585;
wire r6_294;
assign r6_294 = in[5]? r5_588 : r5_587;
wire r6_295;
assign r6_295 = in[5]? r5_590 : r5_589;
wire r6_296;
assign r6_296 = in[5]? r5_592 : r5_591;
wire r6_297;
assign r6_297 = in[5]? r5_594 : r5_593;
wire r6_298;
assign r6_298 = in[5]? r5_596 : r5_595;
wire r6_299;
assign r6_299 = in[5]? r5_598 : r5_597;
wire r6_300;
assign r6_300 = in[5]? r5_600 : r5_599;
wire r6_301;
assign r6_301 = in[5]? r5_602 : r5_601;
wire r6_302;
assign r6_302 = in[5]? r5_604 : r5_603;
wire r6_303;
assign r6_303 = in[5]? r5_606 : r5_605;
wire r6_304;
assign r6_304 = in[5]? r5_608 : r5_607;
wire r6_305;
assign r6_305 = in[5]? r5_610 : r5_609;
wire r6_306;
assign r6_306 = in[5]? r5_612 : r5_611;
wire r6_307;
assign r6_307 = in[5]? r5_614 : r5_613;
wire r6_308;
assign r6_308 = in[5]? r5_616 : r5_615;
wire r6_309;
assign r6_309 = in[5]? r5_618 : r5_617;
wire r6_310;
assign r6_310 = in[5]? r5_620 : r5_619;
wire r6_311;
assign r6_311 = in[5]? r5_622 : r5_621;
wire r6_312;
assign r6_312 = in[5]? r5_624 : r5_623;
wire r6_313;
assign r6_313 = in[5]? r5_626 : r5_625;
wire r6_314;
assign r6_314 = in[5]? r5_628 : r5_627;
wire r6_315;
assign r6_315 = in[5]? r5_630 : r5_629;
wire r6_316;
assign r6_316 = in[5]? r5_632 : r5_631;
wire r6_317;
assign r6_317 = in[5]? r5_634 : r5_633;
wire r6_318;
assign r6_318 = in[5]? r5_636 : r5_635;
wire r6_319;
assign r6_319 = in[5]? r5_638 : r5_637;
wire r6_320;
assign r6_320 = in[5]? r5_640 : r5_639;
wire r6_321;
assign r6_321 = in[5]? r5_642 : r5_641;
wire r7_1;
assign r7_1 = in[6]? r6_2 : r6_1;
wire r7_2;
assign r7_2 = in[6]? r6_4 : r6_3;
wire r7_3;
assign r7_3 = in[6]? r6_6 : r6_5;
wire r7_4;
assign r7_4 = in[6]? r6_8 : r6_7;
wire r7_5;
assign r7_5 = in[6]? r6_10 : r6_9;
wire r7_6;
assign r7_6 = in[6]? r6_12 : r6_11;
wire r7_7;
assign r7_7 = in[6]? r6_14 : r6_13;
wire r7_8;
assign r7_8 = in[6]? r6_16 : r6_15;
wire r7_9;
assign r7_9 = in[6]? r6_18 : r6_17;
wire r7_10;
assign r7_10 = in[6]? r6_20 : r6_19;
wire r7_11;
assign r7_11 = in[6]? r6_22 : r6_21;
wire r7_12;
assign r7_12 = in[6]? r6_24 : r6_23;
wire r7_13;
assign r7_13 = in[6]? r6_26 : r6_25;
wire r7_14;
assign r7_14 = in[6]? r6_28 : r6_27;
wire r7_15;
assign r7_15 = in[6]? r6_30 : r6_29;
wire r7_16;
assign r7_16 = in[6]? r6_32 : r6_31;
wire r7_17;
assign r7_17 = in[6]? r6_34 : r6_33;
wire r7_18;
assign r7_18 = in[6]? r6_36 : r6_35;
wire r7_19;
assign r7_19 = in[6]? r6_38 : r6_37;
wire r7_20;
assign r7_20 = in[6]? r6_40 : r6_39;
wire r7_21;
assign r7_21 = in[6]? r6_42 : r6_41;
wire r7_22;
assign r7_22 = in[6]? r6_44 : r6_43;
wire r7_23;
assign r7_23 = in[6]? r6_46 : r6_45;
wire r7_24;
assign r7_24 = in[6]? r6_48 : r6_47;
wire r7_25;
assign r7_25 = in[6]? r6_50 : r6_49;
wire r7_26;
assign r7_26 = in[6]? r6_52 : r6_51;
wire r7_27;
assign r7_27 = in[6]? r6_54 : r6_53;
wire r7_28;
assign r7_28 = in[6]? r6_56 : r6_55;
wire r7_29;
assign r7_29 = in[6]? r6_58 : r6_57;
wire r7_30;
assign r7_30 = in[6]? r6_60 : r6_59;
wire r7_31;
assign r7_31 = in[6]? r6_62 : r6_61;
wire r7_32;
assign r7_32 = in[6]? r6_64 : r6_63;
wire r7_33;
assign r7_33 = in[6]? r6_66 : r6_65;
wire r7_34;
assign r7_34 = in[6]? r6_68 : r6_67;
wire r7_35;
assign r7_35 = in[6]? r6_70 : r6_69;
wire r7_36;
assign r7_36 = in[6]? r6_72 : r6_71;
wire r7_37;
assign r7_37 = in[6]? r6_74 : r6_73;
wire r7_38;
assign r7_38 = in[6]? r6_76 : r6_75;
wire r7_39;
assign r7_39 = in[6]? r6_78 : r6_77;
wire r7_40;
assign r7_40 = in[6]? r6_80 : r6_79;
wire r7_41;
assign r7_41 = in[6]? r6_82 : r6_81;
wire r7_42;
assign r7_42 = in[6]? r6_84 : r6_83;
wire r7_43;
assign r7_43 = in[6]? r6_86 : r6_85;
wire r7_44;
assign r7_44 = in[6]? r6_88 : r6_87;
wire r7_45;
assign r7_45 = in[6]? r6_90 : r6_89;
wire r7_46;
assign r7_46 = in[6]? r6_92 : r6_91;
wire r7_47;
assign r7_47 = in[6]? r6_94 : r6_93;
wire r7_48;
assign r7_48 = in[6]? r6_96 : r6_95;
wire r7_49;
assign r7_49 = in[6]? r6_98 : r6_97;
wire r7_50;
assign r7_50 = in[6]? r6_100 : r6_99;
wire r7_51;
assign r7_51 = in[6]? r6_102 : r6_101;
wire r7_52;
assign r7_52 = in[6]? r6_104 : r6_103;
wire r7_53;
assign r7_53 = in[6]? r6_106 : r6_105;
wire r7_54;
assign r7_54 = in[6]? r6_108 : r6_107;
wire r7_55;
assign r7_55 = in[6]? r6_110 : r6_109;
wire r7_56;
assign r7_56 = in[6]? r6_112 : r6_111;
wire r7_57;
assign r7_57 = in[6]? r6_114 : r6_113;
wire r7_58;
assign r7_58 = in[6]? r6_116 : r6_115;
wire r7_59;
assign r7_59 = in[6]? r6_118 : r6_117;
wire r7_60;
assign r7_60 = in[6]? r6_120 : r6_119;
wire r7_61;
assign r7_61 = in[6]? r6_122 : r6_121;
wire r7_62;
assign r7_62 = in[6]? r6_124 : r6_123;
wire r7_63;
assign r7_63 = in[6]? r6_126 : r6_125;
wire r7_64;
assign r7_64 = in[6]? r6_128 : r6_127;
wire r7_65;
assign r7_65 = in[6]? r6_130 : r6_129;
wire r7_66;
assign r7_66 = in[6]? r6_132 : r6_131;
wire r7_67;
assign r7_67 = in[6]? r6_134 : r6_133;
wire r7_68;
assign r7_68 = in[6]? r6_136 : r6_135;
wire r7_69;
assign r7_69 = in[6]? r6_138 : r6_137;
wire r7_70;
assign r7_70 = in[6]? r6_140 : r6_139;
wire r7_71;
assign r7_71 = in[6]? r6_142 : r6_141;
wire r7_72;
assign r7_72 = in[6]? r6_144 : r6_143;
wire r7_73;
assign r7_73 = in[6]? r6_146 : r6_145;
wire r7_74;
assign r7_74 = in[6]? r6_148 : r6_147;
wire r7_75;
assign r7_75 = in[6]? r6_150 : r6_149;
wire r7_76;
assign r7_76 = in[6]? r6_152 : r6_151;
wire r7_77;
assign r7_77 = in[6]? r6_154 : r6_153;
wire r7_78;
assign r7_78 = in[6]? r6_156 : r6_155;
wire r7_79;
assign r7_79 = in[6]? r6_158 : r6_157;
wire r7_80;
assign r7_80 = in[6]? r6_160 : r6_159;
wire r7_81;
assign r7_81 = in[6]? r6_162 : r6_161;
wire r7_82;
assign r7_82 = in[6]? r6_164 : r6_163;
wire r7_83;
assign r7_83 = in[6]? r6_166 : r6_165;
wire r7_84;
assign r7_84 = in[6]? r6_168 : r6_167;
wire r7_85;
assign r7_85 = in[6]? r6_170 : r6_169;
wire r7_86;
assign r7_86 = in[6]? r6_172 : r6_171;
wire r7_87;
assign r7_87 = in[6]? r6_174 : r6_173;
wire r7_88;
assign r7_88 = in[6]? r6_176 : r6_175;
wire r7_89;
assign r7_89 = in[6]? r6_178 : r6_177;
wire r7_90;
assign r7_90 = in[6]? r6_180 : r6_179;
wire r7_91;
assign r7_91 = in[6]? r6_182 : r6_181;
wire r7_92;
assign r7_92 = in[6]? r6_184 : r6_183;
wire r7_93;
assign r7_93 = in[6]? r6_186 : r6_185;
wire r7_94;
assign r7_94 = in[6]? r6_188 : r6_187;
wire r7_95;
assign r7_95 = in[6]? r6_190 : r6_189;
wire r7_96;
assign r7_96 = in[6]? r6_192 : r6_191;
wire r7_97;
assign r7_97 = in[6]? r6_194 : r6_193;
wire r7_98;
assign r7_98 = in[6]? r6_196 : r6_195;
wire r7_99;
assign r7_99 = in[6]? r6_198 : r6_197;
wire r7_100;
assign r7_100 = in[6]? r6_200 : r6_199;
wire r7_101;
assign r7_101 = in[6]? r6_202 : r6_201;
wire r7_102;
assign r7_102 = in[6]? r6_204 : r6_203;
wire r7_103;
assign r7_103 = in[6]? r6_206 : r6_205;
wire r7_104;
assign r7_104 = in[6]? r6_208 : r6_207;
wire r7_105;
assign r7_105 = in[6]? r6_210 : r6_209;
wire r7_106;
assign r7_106 = in[6]? r6_212 : r6_211;
wire r7_107;
assign r7_107 = in[6]? r6_214 : r6_213;
wire r7_108;
assign r7_108 = in[6]? r6_216 : r6_215;
wire r7_109;
assign r7_109 = in[6]? r6_218 : r6_217;
wire r7_110;
assign r7_110 = in[6]? r6_220 : r6_219;
wire r7_111;
assign r7_111 = in[6]? r6_222 : r6_221;
wire r7_112;
assign r7_112 = in[6]? r6_224 : r6_223;
wire r7_113;
assign r7_113 = in[6]? r6_226 : r6_225;
wire r7_114;
assign r7_114 = in[6]? r6_228 : r6_227;
wire r7_115;
assign r7_115 = in[6]? r6_230 : r6_229;
wire r7_116;
assign r7_116 = in[6]? r6_232 : r6_231;
wire r7_117;
assign r7_117 = in[6]? r6_234 : r6_233;
wire r7_118;
assign r7_118 = in[6]? r6_236 : r6_235;
wire r7_119;
assign r7_119 = in[6]? r6_238 : r6_237;
wire r7_120;
assign r7_120 = in[6]? r6_240 : r6_239;
wire r7_121;
assign r7_121 = in[6]? r6_242 : r6_241;
wire r7_122;
assign r7_122 = in[6]? r6_244 : r6_243;
wire r7_123;
assign r7_123 = in[6]? r6_246 : r6_245;
wire r7_124;
assign r7_124 = in[6]? r6_248 : r6_247;
wire r7_125;
assign r7_125 = in[6]? r6_250 : r6_249;
wire r7_126;
assign r7_126 = in[6]? r6_252 : r6_251;
wire r7_127;
assign r7_127 = in[6]? r6_254 : r6_253;
wire r7_128;
assign r7_128 = in[6]? r6_256 : r6_255;
wire r7_129;
assign r7_129 = in[6]? r6_258 : r6_257;
wire r7_130;
assign r7_130 = in[6]? r6_260 : r6_259;
wire r7_131;
assign r7_131 = in[6]? r6_262 : r6_261;
wire r7_132;
assign r7_132 = in[6]? r6_264 : r6_263;
wire r7_133;
assign r7_133 = in[6]? r6_266 : r6_265;
wire r7_134;
assign r7_134 = in[6]? r6_268 : r6_267;
wire r7_135;
assign r7_135 = in[6]? r6_270 : r6_269;
wire r7_136;
assign r7_136 = in[6]? r6_272 : r6_271;
wire r7_137;
assign r7_137 = in[6]? r6_274 : r6_273;
wire r7_138;
assign r7_138 = in[6]? r6_276 : r6_275;
wire r7_139;
assign r7_139 = in[6]? r6_278 : r6_277;
wire r7_140;
assign r7_140 = in[6]? r6_280 : r6_279;
wire r7_141;
assign r7_141 = in[6]? r6_282 : r6_281;
wire r7_142;
assign r7_142 = in[6]? r6_284 : r6_283;
wire r7_143;
assign r7_143 = in[6]? r6_286 : r6_285;
wire r7_144;
assign r7_144 = in[6]? r6_288 : r6_287;
wire r7_145;
assign r7_145 = in[6]? r6_290 : r6_289;
wire r7_146;
assign r7_146 = in[6]? r6_292 : r6_291;
wire r7_147;
assign r7_147 = in[6]? r6_294 : r6_293;
wire r7_148;
assign r7_148 = in[6]? r6_296 : r6_295;
wire r7_149;
assign r7_149 = in[6]? r6_298 : r6_297;
wire r7_150;
assign r7_150 = in[6]? r6_300 : r6_299;
wire r7_151;
assign r7_151 = in[6]? r6_302 : r6_301;
wire r7_152;
assign r7_152 = in[6]? r6_304 : r6_303;
wire r7_153;
assign r7_153 = in[6]? r6_306 : r6_305;
wire r7_154;
assign r7_154 = in[6]? r6_308 : r6_307;
wire r7_155;
assign r7_155 = in[6]? r6_310 : r6_309;
wire r7_156;
assign r7_156 = in[6]? r6_312 : r6_311;
wire r7_157;
assign r7_157 = in[6]? r6_314 : r6_313;
wire r7_158;
assign r7_158 = in[6]? r6_316 : r6_315;
wire r7_159;
assign r7_159 = in[6]? r6_318 : r6_317;
wire r7_160;
assign r7_160 = in[6]? r6_320 : r6_319;
assign r7_161 = r6_321;
wire r8_1;
assign r8_1 = in[7]? r7_2 : r7_1;
wire r8_2;
assign r8_2 = in[7]? r7_4 : r7_3;
wire r8_3;
assign r8_3 = in[7]? r7_6 : r7_5;
wire r8_4;
assign r8_4 = in[7]? r7_8 : r7_7;
wire r8_5;
assign r8_5 = in[7]? r7_10 : r7_9;
wire r8_6;
assign r8_6 = in[7]? r7_12 : r7_11;
wire r8_7;
assign r8_7 = in[7]? r7_14 : r7_13;
wire r8_8;
assign r8_8 = in[7]? r7_16 : r7_15;
wire r8_9;
assign r8_9 = in[7]? r7_18 : r7_17;
wire r8_10;
assign r8_10 = in[7]? r7_20 : r7_19;
wire r8_11;
assign r8_11 = in[7]? r7_22 : r7_21;
wire r8_12;
assign r8_12 = in[7]? r7_24 : r7_23;
wire r8_13;
assign r8_13 = in[7]? r7_26 : r7_25;
wire r8_14;
assign r8_14 = in[7]? r7_28 : r7_27;
wire r8_15;
assign r8_15 = in[7]? r7_30 : r7_29;
wire r8_16;
assign r8_16 = in[7]? r7_32 : r7_31;
wire r8_17;
assign r8_17 = in[7]? r7_34 : r7_33;
wire r8_18;
assign r8_18 = in[7]? r7_36 : r7_35;
wire r8_19;
assign r8_19 = in[7]? r7_38 : r7_37;
wire r8_20;
assign r8_20 = in[7]? r7_40 : r7_39;
wire r8_21;
assign r8_21 = in[7]? r7_42 : r7_41;
wire r8_22;
assign r8_22 = in[7]? r7_44 : r7_43;
wire r8_23;
assign r8_23 = in[7]? r7_46 : r7_45;
wire r8_24;
assign r8_24 = in[7]? r7_48 : r7_47;
wire r8_25;
assign r8_25 = in[7]? r7_50 : r7_49;
wire r8_26;
assign r8_26 = in[7]? r7_52 : r7_51;
wire r8_27;
assign r8_27 = in[7]? r7_54 : r7_53;
wire r8_28;
assign r8_28 = in[7]? r7_56 : r7_55;
wire r8_29;
assign r8_29 = in[7]? r7_58 : r7_57;
wire r8_30;
assign r8_30 = in[7]? r7_60 : r7_59;
wire r8_31;
assign r8_31 = in[7]? r7_62 : r7_61;
wire r8_32;
assign r8_32 = in[7]? r7_64 : r7_63;
wire r8_33;
assign r8_33 = in[7]? r7_66 : r7_65;
wire r8_34;
assign r8_34 = in[7]? r7_68 : r7_67;
wire r8_35;
assign r8_35 = in[7]? r7_70 : r7_69;
wire r8_36;
assign r8_36 = in[7]? r7_72 : r7_71;
wire r8_37;
assign r8_37 = in[7]? r7_74 : r7_73;
wire r8_38;
assign r8_38 = in[7]? r7_76 : r7_75;
wire r8_39;
assign r8_39 = in[7]? r7_78 : r7_77;
wire r8_40;
assign r8_40 = in[7]? r7_80 : r7_79;
wire r8_41;
assign r8_41 = in[7]? r7_82 : r7_81;
wire r8_42;
assign r8_42 = in[7]? r7_84 : r7_83;
wire r8_43;
assign r8_43 = in[7]? r7_86 : r7_85;
wire r8_44;
assign r8_44 = in[7]? r7_88 : r7_87;
wire r8_45;
assign r8_45 = in[7]? r7_90 : r7_89;
wire r8_46;
assign r8_46 = in[7]? r7_92 : r7_91;
wire r8_47;
assign r8_47 = in[7]? r7_94 : r7_93;
wire r8_48;
assign r8_48 = in[7]? r7_96 : r7_95;
wire r8_49;
assign r8_49 = in[7]? r7_98 : r7_97;
wire r8_50;
assign r8_50 = in[7]? r7_100 : r7_99;
wire r8_51;
assign r8_51 = in[7]? r7_102 : r7_101;
wire r8_52;
assign r8_52 = in[7]? r7_104 : r7_103;
wire r8_53;
assign r8_53 = in[7]? r7_106 : r7_105;
wire r8_54;
assign r8_54 = in[7]? r7_108 : r7_107;
wire r8_55;
assign r8_55 = in[7]? r7_110 : r7_109;
wire r8_56;
assign r8_56 = in[7]? r7_112 : r7_111;
wire r8_57;
assign r8_57 = in[7]? r7_114 : r7_113;
wire r8_58;
assign r8_58 = in[7]? r7_116 : r7_115;
wire r8_59;
assign r8_59 = in[7]? r7_118 : r7_117;
wire r8_60;
assign r8_60 = in[7]? r7_120 : r7_119;
wire r8_61;
assign r8_61 = in[7]? r7_122 : r7_121;
wire r8_62;
assign r8_62 = in[7]? r7_124 : r7_123;
wire r8_63;
assign r8_63 = in[7]? r7_126 : r7_125;
wire r8_64;
assign r8_64 = in[7]? r7_128 : r7_127;
wire r8_65;
assign r8_65 = in[7]? r7_130 : r7_129;
wire r8_66;
assign r8_66 = in[7]? r7_132 : r7_131;
wire r8_67;
assign r8_67 = in[7]? r7_134 : r7_133;
wire r8_68;
assign r8_68 = in[7]? r7_136 : r7_135;
wire r8_69;
assign r8_69 = in[7]? r7_138 : r7_137;
wire r8_70;
assign r8_70 = in[7]? r7_140 : r7_139;
wire r8_71;
assign r8_71 = in[7]? r7_142 : r7_141;
wire r8_72;
assign r8_72 = in[7]? r7_144 : r7_143;
wire r8_73;
assign r8_73 = in[7]? r7_146 : r7_145;
wire r8_74;
assign r8_74 = in[7]? r7_148 : r7_147;
wire r8_75;
assign r8_75 = in[7]? r7_150 : r7_149;
wire r8_76;
assign r8_76 = in[7]? r7_152 : r7_151;
wire r8_77;
assign r8_77 = in[7]? r7_154 : r7_153;
wire r8_78;
assign r8_78 = in[7]? r7_156 : r7_155;
wire r8_79;
assign r8_79 = in[7]? r7_158 : r7_157;
wire r8_80;
assign r8_80 = in[7]? r7_160 : r7_159;
assign r8_81 = r6_161;
wire r9_1;
assign r9_1 = in[8]? r8_2 : r8_1;
wire r9_2;
assign r9_2 = in[8]? r8_4 : r8_3;
wire r9_3;
assign r9_3 = in[8]? r8_6 : r8_5;
wire r9_4;
assign r9_4 = in[8]? r8_8 : r8_7;
wire r9_5;
assign r9_5 = in[8]? r8_10 : r8_9;
wire r9_6;
assign r9_6 = in[8]? r8_12 : r8_11;
wire r9_7;
assign r9_7 = in[8]? r8_14 : r8_13;
wire r9_8;
assign r9_8 = in[8]? r8_16 : r8_15;
wire r9_9;
assign r9_9 = in[8]? r8_18 : r8_17;
wire r9_10;
assign r9_10 = in[8]? r8_20 : r8_19;
wire r9_11;
assign r9_11 = in[8]? r8_22 : r8_21;
wire r9_12;
assign r9_12 = in[8]? r8_24 : r8_23;
wire r9_13;
assign r9_13 = in[8]? r8_26 : r8_25;
wire r9_14;
assign r9_14 = in[8]? r8_28 : r8_27;
wire r9_15;
assign r9_15 = in[8]? r8_30 : r8_29;
wire r9_16;
assign r9_16 = in[8]? r8_32 : r8_31;
wire r9_17;
assign r9_17 = in[8]? r8_34 : r8_33;
wire r9_18;
assign r9_18 = in[8]? r8_36 : r8_35;
wire r9_19;
assign r9_19 = in[8]? r8_38 : r8_37;
wire r9_20;
assign r9_20 = in[8]? r8_40 : r8_39;
assign r9_21 = r8_41;
wire r10_1;
assign r10_1 = in[9]? r9_2 : r9_1;
wire r10_2;
assign r10_2 = in[9]? r9_4 : r9_3;
wire r10_3;
assign r10_3 = in[9]? r9_6 : r9_5;
wire r10_4;
assign r10_4 = in[9]? r9_8 : r9_7;
wire r10_5;
assign r10_5 = in[9]? r9_10 : r9_9;
wire r10_6;
assign r10_6 = in[9]? r9_12 : r9_11;
wire r10_7;
assign r10_7 = in[9]? r9_14 : r9_13;
wire r10_8;
assign r10_8 = in[9]? r9_16 : r9_15;
wire r10_9;
assign r10_9 = in[9]? r9_18 : r9_17;
wire r10_10;
assign r10_10 = in[9]? r9_20 : r9_19;
assign r10_11 = r9_21;
wire r11_1;
assign r11_1 = in[10]? r10_2 : r10_1;
wire r11_2;
assign r11_2 = in[10]? r10_4 : r10_3;
wire r11_3;
assign r11_3 = in[10]? r10_6 : r10_5;
wire r11_4;
assign r11_4 = in[10]? r10_8 : r10_7;
wire r11_5;
assign r11_5 = in[10]? r10_10 : r10_9;
assign r11_6 = r10_11;
wire r12_1;
assign r12_1 = in[11]? r11_2 : r11_1;
wire r12_2;
assign r12_2 = in[11]? r11_4 : r11_3;
wire r12_3;
assign r12_3 = in[11]? r11_6 : r11_5;
wire r13_1;
assign r13_1 = in[12]? r12_2 : r12_1;
assign r13_2 = r12_3;
wire r;
assign r = in[13]? r13_2 : r13_1;

endmodule
