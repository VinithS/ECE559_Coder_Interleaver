`timescale 1ns / 1ps

module coder_interleaver_tb();

	//instantiate modules
	reg size_6144, clk, rst, shift_en, ready_in;
	reg [6143:0] input_val;
	wire [6143:0] out_val;
	
	reg [7:0] byte_in;
//11011111
	wire outi, outpii;
	//monitor output i

	interleaver_top_level_early_test inter_inst(
	.k_size_6144(size_6144),      // 0 if 1056, 1 if 6144 block size
	.databyte_in(byte_in),  // byte-wise serial input
	.clock(clk),         // clock 
	.rst(rst),			// reset
	.shift_en(shift_en),
	.ready_in(ready_in),       // asserted to indicate the whole block is filled and this module starts output serial stream; as of now it needs to be asserted for at least K cycles
	.outi(outi), // bitserial output using the same sequence as input, i.e. ci
	.outpii(outpii) // bitserial output after remapping, i.e. cpii
	//output process_complete
	);
	
	//assert inside wires potentially interested in
	wire [6151:0] p_shift_reg_out;
	assign p_shift_reg_out = inter_inst.shift_reg_out;
	wire [6143:0] p_reg_buf_out;
	assign  p_reg_buf_out= inter_inst.reg_buf_out;

	wire [6143:0] p_ci_array, p_cpii_array;
	assign  p_ci_array= inter_inst.ci_array;
	assign  p_cpii_array= inter_inst.cpii_array;

	wire [13:0] mux_ind;
	assign mux_ind = inter_inst.mux_ind;
integer i = 0;
	initial begin
		clk=0;
		rst=0;
		byte_in=8'b11011111;
		shift_en=0;
		ready_in=0;
		size_6144=1;
		@(negedge clk);
		rst=1;
		@(negedge clk);
		rst=0;

		//start shifting in
		@(negedge clk);
		shift_en=1;
		for (i=0; i < 769; i=i+1) begin
			@(negedge clk) $display("shifting cycle: %d",i);
		end
		shift_en=0;
		$display("finished shifting");
		//want to check the input and output now
		$display("shiftregister output is %b",p_shift_reg_out);

		@(negedge clk) ready_in=1;
		$display("time%d, ready_in asserted",$time);
		@(negedge clk) ready_in=0;
		@(negedge clk) ready_in=0;
		@(negedge clk) ready_in=0;
		$display("secondary buffer output is %b",p_reg_buf_out);
		
		$display("ciarray is %b",p_ci_array);
		$display("cpiiarray is %b",p_cpii_array);
		$stop;
		for (i = 0; i < 6144; i=i+1) begin
			@(negedge clk) $display("ready_in cycle: %d",i);
			$display("Time:%d, mux index:%d, \t Outi %b,\tOutPii: %b",$time,mux_ind, outi,outpii);
		end
		//shifting now
		//interested in mux_ind
		#1000; // wait 50 ns
		// input_val = 6144'b110110011000001110010010101011111001000001010010110111001110110010111010000000111001101110100010001010101111110001111000011100100111101011100111110011100000101011010101010110100000000000100111011100000000010100110001110011100101111011101000001011111000111001001101110011000111001010011111101110001011110100010110000011010111101010000001000100100000011110010001100011100111101010000000000001101101010010010111011000000111101110100000011000100010110001101111101110010001011110111100010010001101000001100101101010110011101000101111111010100110111011000110100000101010100000111010111011100100111110110001001100110010001110011011111111110011101010000101110101100001110100101111001010100010101001101110011001101000010110011101100010110100110101001100010001001010001111100100001100001111010001011010111101011000011100110000001011100001011010101001001100111001100010110010001111101010111111011100010101010010100010110010110010001110000100011110101101011111011001001110101111001101000110100101100011010011010001110000111011111100000010010011101101101010110001110100110110100011111110110100101001010010010101100110001010110011001111110100111101000001001010010111000001110101001010111001011111001001111100101010001101111011111000101010101100100001110000101110001001111011100010011111110100110010000010111000000011110011111100001010101011001110001100100001111001000111010000000101111111110111001110001001011001100110001110100101000000010011000000011010110010000010000000101111100010001100110110100111111011110101100001011101100111011100011011110001011111101001011101101001101010010111000011001001111110000001011101000010100010001110111111010110111000001100000110110101110100110010110000110001001001110111001011000111010101100100101101100101010011010011000100011101010000110000100000000100110101000010101000101100100010100001011100111011001101110010111101011111000011001011000100010001100101001110110101111011001001100100110100100000001100110001010011001001111101101100111010010110101111001101011101010100010100111110111100110010010011001010000100100010001110010001110101010011011100010100110001100001001100011111110100110101000110001101110000010001110100111000101001000000001111101111100101000000111010100001010100011010110010111111010100011101101011110111101010101011101100010101000100111101001111010011111100011010010111011100101010100110100011000101000111101101011000001000000000001110110101011000111101110000011010111111111000110100100100101100001101101101001100101111101011101110011011000001101111110011010000101010001011001101011001001001110101001001010011111000011100110111110101100100110010011001000000010111100011111011110100011001101100111001011101011110001001000111011011010010111101111001011110000110000001001101100010110000010110111101011111001111111000011001111100110100110100100110000010100111111011100110010011101010111001011010100101101001100001001111011101000001000101000101101110001101010001010000110011000110100111000010110111111011000111010011100001111100010011101000001111111110011000100011011111000110001111111101011100111011111010111011110111010110001011100010100101101011000000101110010010011100101111011001101011011110101101001000001010100011111101110010011001000000100001111101000000010111011110010100101001100101001101111001101010001100100011100001001011001100001010000000101101000100110111111001000001011111110001100101011101100111011010010110111000010110111110010011001010011110001010101011101011001110101011011111111000101110001001101001011000111001110100000001010000110111110100111110100010111010010010011000111010110100011111000100001010100100000100111001110101111111111101110110111101010001100101111100110011010110000010101110000010101100010100111000010011011010100111101110010001011011111010100111000011101000111111001111111010101010011000010011000101101000101010101101000011010111010001111010110101110110001010010110000100001110000001001110011011110011001000100011011001001110000110001111101100011111001101001010111011001011111101000000001001101001101000010001110100111010010011000110000011101010111101111010110000001001111001100011111000101011100001011100111100100001111111111111011110100011101001101101100011110001101111100100000010110111011001001001100101001111001100000010001100001001000110110010000000100111000000110011011000011101101010001100010011010000111110011111101010100001001001100101000011100110000111011101011101010010001011010111010000101111000010100110110101011111101101010000001011100111010001010011110001100000101010000100000101001001001001101011110100010001110111001011000111010110111011000100101111010001001101101010100011011000011100110101001010111011100110100011101010000010010110011111111111010100001011100101101001001011110101100100001110111101001001100010101101011011101111011100100111110110001001011001001011000100111000110100010001100001101001100000100110110010000110010111111101001101111100000110011000110110110100001000000110011010111001100110100010100111010011011111111010111100110101111010011010011111000100110101101111011100010011011010000101111111101100011010100010110011000101000101100010101101000110101011100010111111011111000101111101011110101101000010000100000110000001100001010011001000000001111000001010000111001110010000001111100110010001101010111000001111000010110000010011101111101111000011101100110000010011011010110100010110000001010010101000010111010101110010110010001000000110110011001101000101110111000111101001000110101001110001111011100001011100000100111100100010111111111011001110100010001110111110111001011010001010001010111010110110101110101100010101001101000000100011011101000010010011011001100000000001000100100100100110110110010011111010010001101001010101001000010110011000111010111000111010101011111100100110100000100011101110100001111001010100000101000110001110000110001110101100011011100010011011110001011001101010110101011100001101100100000100111011110010000000100101101101100110101111001001001101110011011111001111111100000001101110101110001111101011011111101010101001010100111011000000011000101100010000001111101100001100111111000001010110111001100000010100110111000100000000001000110001110111001000010011100001111000101001001010101110010100000011100111011110; // 0000..<6136> more zeros..0001
		// size_6144 = 1;
		// theoretic out: 011100100000011101110011010100111101010000101000001000111011101111111100011110011100100000101111011010011001100100001100010000011101011110110011111000111010001010000011100111000010100010000100011000010010110111010110110011100000011011111000011011010011000001111001101011110010000111000011100111110111101001110001000110000000100110011000101011001010100111000001011011011110101000110000111010000111111001100110010001100001010001111010100101011011001110110110101000001001100100011001000010010000111011011111110001001100100110011011101110110010011101100001111101010100000110011111110100101000010101110011101000011111001000101101001000110001100001001101010001001010000111110001001110111000111111011000100110001100011110011010010101000100010100000001010011111001010110001011010001001100111000111111100101011101110010100100010111010010000101010000111010110100000010100111010100111111100111100100110000110011101010100101001101101110101000110111001100111100011101100001110111111100010001011111111000110101000111001010000010011100001101101100100100011001111101001010000111110010011101011110000011011100101101011101000111110100100111100100000100101000000101010101001100110010111011011011100101000101001111010100101001010011011011001000111010100110101000110000000110110011101000011101110110111010110011001100000110011001111000101111101011001110100101111111111111000011000110011111111010111100100000111010100101000000000101011101001100000001010100110000010101100111011011110011011111010110101001000010100110010110101101000000110010110011101000001011111011000011001010001100101100110111001011101101010101010011000010100010111101101101100100110000000100010111000100011010010100101101010111111101100110011011101100011100100011111010110110110001111100100110011001010110001111100111010100000000010100010111111000001010100101110001101010011011010011100011101101101101011000001111001000000101010110000110110011000010011110011000110000110110001100100001110001111101100001111111101010010000101010001000101100110100110000111100101001001101110100111100011000111000001000111011001000001101101100010001011111010000001110100100000011101101010110100011000110100000101110011011001110001101100000011100010011110010000101100010100010011000011000110011111100100000011000000111100101110011111111010110110111011010001000010000111110101100010110100100010101001000111100111001100100110101011011101011010010010000010010110111001111111000001110110101110111110100110101001010001101101110010100110000111111100110001010100001010100111100010011011001100101111110010111000001100110000010110011000011000010110000100100011001000110110011111111000011111110011111011101001111111111101101100100011001010011001011101110011111100111111111010001000000100110110011000110001101010011001000010111101001000001111000101101010101001100000110101000111101111111001011111100000011111010000111111010101110010101001100101111100001011101100111000111001101100110011111110111111000100001011101011100010010111001011110110000000011100110010010100001110010001110110101100000010011111110100000100101111100001011111011111111110111111110111001011101100100000110011011001101111101010110000100110100111001100110010101110011001010000110100100011111100010000010101110101001000110010100110011111101000111000101100100101010101111110001010100111110100000000111001000101010001000000010111111101100100100111101100100010001101000001110001110000101101110011000101011000000001101101101110110110100000010100100011010001111011100001011101000001001000110000101100001110011101101000000000000011010100101111010010101010100111111001011100010100000010110111010010101001101001101101111010110000010110101100010010111110011110001101001000010011001100100110111100110001010100101110010001000011010100011010100110100000111110011100011111001101110011000100110100110100000001010011001100010111010001011110101011011001101000011011101011010001001101000000101101000000100001001010000011110011000110001111010000000110000010010101000111011010100100111001111110011101001011000001010100101000101001110011100000110100001000111110010011010101111010110111101111011010100100111000000111011010100110101110111011000011010100111001011100001111100110101010101011111100001000110011010001000110001010001100100000000001111100111011000000011101110010011110100010011110011111010000011100000000100101101111000011011101110111111110101011100010001101001110000001011000001111011010001101111100101010101100000100010000001010010101110111001110101100001101010111101101001111101000001010101011011111001010110111011101011100101010000000101010010000011000111001111000100010000101000100110011000100000000111101110001101001111110000010011100000110011000001100110100101100001111101010110010101000111010101011000100111011000010110010001001101011011000000100001111111101111111111001101010101101011110000011100101111100101010011100101100101101000101001011010000000001111100010010100011011000101101110011000100010110100101001101101101011110001110001110011011111011001111100100101101011100111111110010001100111110100000011101011001000101100000000011111101100100111111111110011111001110011111000011010110010010111100101000111011111101010000001101001011111110100110010010101010010001000000100010111011001010111110010100100011000100011010000011100100001110111111011101101011101001110111110100010011101010100000111001111111101110001101110011010110111110111111100011010100001001110011001100110100101010001100010010100111000010010000100001010001110101100111100110010110110001110000101100111001011111110000010001101000111101011000100010101010011110000001000100100110011111010011001110110001100101001011010000001011001101100011100001000011110111101110011001101010001100111010110111001000111101110011110110110011011111011010101110101111110011000011000010010101001000001100111110110111101000101110100001001110000010001100110100100100010000001100100101111100000001101101011110011001111111101011001111100011001010110111011110101101100011111010100110110100101111001011110011111111100000011000100101000100001010110111001010010110110110111100011110011000001100000101010101010110111001010100010010011111000111100111100111001101001011010000111100010101000000011011011011111111101100101010110001101
		// 60 output bits: 101100011010101001101111111110110110110000000101010001111000...
		// Matches the output last 60 bits of the python script.
		

		// #1000; // wait 50 ns
		// input_val = 1056'b010111110010101000110110111010010001110100001010001001010011110001101111001001110010110100111100000010111001011111010100000000000001101001110100000010100111100111111110001101100110101011111111110011000111011010111100101000100110000001000000011101000110100100001010010001100000100010111100001010011000011100111011010100110101000000010101110001000001001011110111001101110001010100010100000010111101011001000000000100001000011000100100000111010010010000000111011011011011000001110000100010110011100100011010110101100101101110001000111011101111010111010100001111011000010111100100011010011000001110010000001001000011010100000010111101111101110000000110001010011001110010001111001100000010110011111011011010010111000010101101001110010011011010110001111100100000011100101101011001111101111101101110111001001001111110110011110010010110110001001011010100000100011111001000000111000001101111100110011101000010011110111100001011101000011111100011100010001100010010101100100010000111011100100110000101000001010001101011001010110110100110010000011010100100000001100100;
		// size_6144 = 0;
		// theoretic out: 001010100100000111010100000001000010000011111001011110101000111111000001010101000110000011001010000111100100001000001101101010000100001110110001111100111110110100001001100111100100100011101100011011011001001000000011000001110011110001011110011101111010101110110000000011001011000011010010001110000100010011100001001001000001011010101010000110001011000100111011011101001001001001010011011101001011100010010010100000011011000101001100011100010010000100110001101110011001111000001100000101010110011000110111101110110101100001111000000001101110101110001111010100000100100111100010110000101010001010110001111101110010100011001110100100000111111001110000011100101010100000010010101101111001001110001101101001101001111111111110000011101111000110111110001000000110101111111001101100010000100100011100010100010111111001000000011010101100100101110001001111111110011101101001011000101010010010001011111010000101101101110000111101010011101101010001001000000111100000010000010011011010110010110000011101111111000101010000100110010010101011111111001000010101100000100011
		#1000;
	end
	
	/* First test with input value 1 with a large size */
	// initial begin
	// 	// $display("input_val: %b",input_val);
	// 	// $display("\ttime,\tinputval,\tsize_6144,\tout_val");
	// 	// $monitor("Time:%d, Outi %b,\tOutPii: %b",$time,outi,outpii);
	// end
	
//	initial begin
//		$display("\ttime,\tinputval,\tsize_6144,\tout_val");
//		$monitor("%d,\t%h,\t%b,\t%h",$time,input_val, size_6144, out_val);
//	end
	always 
		#5 clk=~clk;


endmodule
