`ifndef CODER_INTERLEAVER_H
`define CODER_INTERLEAVER_H

module coder_interleaver (
	input [6143:0] cin,    // Clock
	input K_eq_6144,
	output [6143:0] cout
);
	
	wire [6143:0] cj_6144, cj_1056;

// module mux2to1 (
// 	input in_a, in_b,    // Clock
// 	input sel, // Clock Enable
// 	input out,  // Asynchronous reset active low
// );

parameter f1_6144=263;

parameter f1_1056=17;

parameter f2_6144=480;

parameter f2_1056=66;





//for j from 0 to 6143
genvar  j;
generate
	for (j=0;j<4800;j=j+1)
	begin: loop0to4799
		assign cout[j]=K_eq_6144?cj_6144[j]:cj_1056[j];
	end
endgenerate

//for j2 from 0 to 6143
genvar  j2;
generate
	for (j2=4800;j2<6144;j2=j2+1)
	begin: loop4800to6143
		assign cout[j2]=K_eq_6144?cj_6144[j2]:cj_1056[j2];
	end
endgenerate

//for j from 0 to 1055

// cj_6144[j]=cin[(f1_6144*j+f2_6144*j*j)%6144]

// cj_1056[j]=cin[(f1_1056*j+f2_1056*j*j)%1056]

genvar  i1;
generate
	for (i1=0;i1<1056;i1=i1+1)
	begin: loop0to1055
		assign cj_6144[i1]=cin[(f1_6144*i1+f2_6144*i1*i1)%6144];
		assign cj_1056[i1]=cin[(f1_1056*i1+f2_1056*i1*i1)%1056];
	end
endgenerate


//for j from 1056 to 6143
genvar  i2;
generate
	for (i2=1056;i2<2100;i2=i2+1)
	begin: loop1056to6143
		assign cj_6144[i2]=cin[(f1_6144*i2+f2_6144*i2*i2)%6144];
		assign cj_1056[i2]=1'b0;
	end
endgenerate

genvar  i3;
generate
	for (i3=2100;i3<6144;i3=i3+1)
	begin: loop1056to6144
		//assign cj_6144[i3]=cin[(f1_6144*i3+f2_6144*i3*i3)%6144];
		assign cj_1056[i3]=1'b0;
	end
endgenerate



assign cj_6144[2100] = cin[876];
assign cj_6144[2101] = cin[2387];
assign cj_6144[2102] = cin[4858];
assign cj_6144[2103] = cin[2145];
assign cj_6144[2104] = cin[392];
assign cj_6144[2105] = cin[5743];
assign cj_6144[2106] = cin[5910];
assign cj_6144[2107] = cin[893];
assign cj_6144[2108] = cin[2980];
assign cj_6144[2109] = cin[6027];
assign cj_6144[2110] = cin[3890];
assign cj_6144[2111] = cin[2713];
assign cj_6144[2112] = cin[2496];
assign cj_6144[2113] = cin[3239];
assign cj_6144[2114] = cin[4942];
assign cj_6144[2115] = cin[1461];
assign cj_6144[2116] = cin[5084];
assign cj_6144[2117] = cin[3523];
assign cj_6144[2118] = cin[2922];
assign cj_6144[2119] = cin[3281];
assign cj_6144[2120] = cin[4600];
assign cj_6144[2121] = cin[735];
assign cj_6144[2122] = cin[3974];
assign cj_6144[2123] = cin[2029];
assign cj_6144[2124] = cin[1044];
assign cj_6144[2125] = cin[1019];
assign cj_6144[2126] = cin[1954];
assign cj_6144[2127] = cin[3849];
assign cj_6144[2128] = cin[560];
assign cj_6144[2129] = cin[4375];
assign cj_6144[2130] = cin[3006];
assign cj_6144[2131] = cin[2597];
assign cj_6144[2132] = cin[3148];
assign cj_6144[2133] = cin[4659];
assign cj_6144[2134] = cin[986];
assign cj_6144[2135] = cin[4417];
assign cj_6144[2136] = cin[2664];
assign cj_6144[2137] = cin[1871];
assign cj_6144[2138] = cin[2038];
assign cj_6144[2139] = cin[3165];
assign cj_6144[2140] = cin[5252];
assign cj_6144[2141] = cin[2155];
assign cj_6144[2142] = cin[18];
assign cj_6144[2143] = cin[4985];
assign cj_6144[2144] = cin[4768];
assign cj_6144[2145] = cin[5511];
assign cj_6144[2146] = cin[1070];
assign cj_6144[2147] = cin[3733];
assign cj_6144[2148] = cin[1212];
assign cj_6144[2149] = cin[5795];
assign cj_6144[2150] = cin[5194];
assign cj_6144[2151] = cin[5553];
assign cj_6144[2152] = cin[728];
assign cj_6144[2153] = cin[3007];
assign cj_6144[2154] = cin[102];
assign cj_6144[2155] = cin[4301];
assign cj_6144[2156] = cin[3316];
assign cj_6144[2157] = cin[3291];
assign cj_6144[2158] = cin[4226];
assign cj_6144[2159] = cin[6121];
assign cj_6144[2160] = cin[2832];
assign cj_6144[2161] = cin[503];
assign cj_6144[2162] = cin[5278];
assign cj_6144[2163] = cin[4869];
assign cj_6144[2164] = cin[5420];
assign cj_6144[2165] = cin[787];
assign cj_6144[2166] = cin[3258];
assign cj_6144[2167] = cin[545];
assign cj_6144[2168] = cin[4936];
assign cj_6144[2169] = cin[4143];
assign cj_6144[2170] = cin[4310];
assign cj_6144[2171] = cin[5437];
assign cj_6144[2172] = cin[1380];
assign cj_6144[2173] = cin[4427];
assign cj_6144[2174] = cin[2290];
assign cj_6144[2175] = cin[1113];
assign cj_6144[2176] = cin[896];
assign cj_6144[2177] = cin[1639];
assign cj_6144[2178] = cin[3342];
assign cj_6144[2179] = cin[6005];
assign cj_6144[2180] = cin[3484];
assign cj_6144[2181] = cin[1923];
assign cj_6144[2182] = cin[1322];
assign cj_6144[2183] = cin[1681];
assign cj_6144[2184] = cin[3000];
assign cj_6144[2185] = cin[5279];
assign cj_6144[2186] = cin[2374];
assign cj_6144[2187] = cin[429];
assign cj_6144[2188] = cin[5588];
assign cj_6144[2189] = cin[5563];
assign cj_6144[2190] = cin[354];
assign cj_6144[2191] = cin[2249];
assign cj_6144[2192] = cin[5104];
assign cj_6144[2193] = cin[2775];
assign cj_6144[2194] = cin[1406];
assign cj_6144[2195] = cin[997];
assign cj_6144[2196] = cin[1548];
assign cj_6144[2197] = cin[3059];
assign cj_6144[2198] = cin[5530];
assign cj_6144[2199] = cin[2817];
assign cj_6144[2200] = cin[1064];
assign cj_6144[2201] = cin[271];
assign cj_6144[2202] = cin[438];
assign cj_6144[2203] = cin[1565];
assign cj_6144[2204] = cin[3652];
assign cj_6144[2205] = cin[555];
assign cj_6144[2206] = cin[4562];
assign cj_6144[2207] = cin[3385];
assign cj_6144[2208] = cin[3168];
assign cj_6144[2209] = cin[3911];
assign cj_6144[2210] = cin[5614];
assign cj_6144[2211] = cin[2133];
assign cj_6144[2212] = cin[5756];
assign cj_6144[2213] = cin[4195];
assign cj_6144[2214] = cin[3594];
assign cj_6144[2215] = cin[3953];
assign cj_6144[2216] = cin[5272];
assign cj_6144[2217] = cin[1407];
assign cj_6144[2218] = cin[4646];
assign cj_6144[2219] = cin[2701];
assign cj_6144[2220] = cin[1716];
assign cj_6144[2221] = cin[1691];
assign cj_6144[2222] = cin[2626];
assign cj_6144[2223] = cin[4521];
assign cj_6144[2224] = cin[1232];
assign cj_6144[2225] = cin[5047];
assign cj_6144[2226] = cin[3678];
assign cj_6144[2227] = cin[3269];
assign cj_6144[2228] = cin[3820];
assign cj_6144[2229] = cin[5331];
assign cj_6144[2230] = cin[1658];
assign cj_6144[2231] = cin[5089];
assign cj_6144[2232] = cin[3336];
assign cj_6144[2233] = cin[2543];
assign cj_6144[2234] = cin[2710];
assign cj_6144[2235] = cin[3837];
assign cj_6144[2236] = cin[5924];
assign cj_6144[2237] = cin[2827];
assign cj_6144[2238] = cin[690];
assign cj_6144[2239] = cin[5657];
assign cj_6144[2240] = cin[5440];
assign cj_6144[2241] = cin[39];
assign cj_6144[2242] = cin[1742];
assign cj_6144[2243] = cin[4405];
assign cj_6144[2244] = cin[1884];
assign cj_6144[2245] = cin[323];
assign cj_6144[2246] = cin[5866];
assign cj_6144[2247] = cin[81];
assign cj_6144[2248] = cin[1400];
assign cj_6144[2249] = cin[3679];
assign cj_6144[2250] = cin[774];
assign cj_6144[2251] = cin[4973];
assign cj_6144[2252] = cin[3988];
assign cj_6144[2253] = cin[3963];
assign cj_6144[2254] = cin[4898];
assign cj_6144[2255] = cin[649];
assign cj_6144[2256] = cin[3504];
assign cj_6144[2257] = cin[1175];
assign cj_6144[2258] = cin[5950];
assign cj_6144[2259] = cin[5541];
assign cj_6144[2260] = cin[6092];
assign cj_6144[2261] = cin[1459];
assign cj_6144[2262] = cin[3930];
assign cj_6144[2263] = cin[1217];
assign cj_6144[2264] = cin[5608];
assign cj_6144[2265] = cin[4815];
assign cj_6144[2266] = cin[4982];
assign cj_6144[2267] = cin[6109];
assign cj_6144[2268] = cin[2052];
assign cj_6144[2269] = cin[5099];
assign cj_6144[2270] = cin[2962];
assign cj_6144[2271] = cin[1785];
assign cj_6144[2272] = cin[1568];
assign cj_6144[2273] = cin[2311];
assign cj_6144[2274] = cin[4014];
assign cj_6144[2275] = cin[533];
assign cj_6144[2276] = cin[4156];
assign cj_6144[2277] = cin[2595];
assign cj_6144[2278] = cin[1994];
assign cj_6144[2279] = cin[2353];
assign cj_6144[2280] = cin[3672];
assign cj_6144[2281] = cin[5951];
assign cj_6144[2282] = cin[3046];
assign cj_6144[2283] = cin[1101];
assign cj_6144[2284] = cin[116];
assign cj_6144[2285] = cin[91];
assign cj_6144[2286] = cin[1026];
assign cj_6144[2287] = cin[2921];
assign cj_6144[2288] = cin[5776];
assign cj_6144[2289] = cin[3447];
assign cj_6144[2290] = cin[2078];
assign cj_6144[2291] = cin[1669];
assign cj_6144[2292] = cin[2220];
assign cj_6144[2293] = cin[3731];
assign cj_6144[2294] = cin[58];
assign cj_6144[2295] = cin[3489];
assign cj_6144[2296] = cin[1736];
assign cj_6144[2297] = cin[943];
assign cj_6144[2298] = cin[1110];
assign cj_6144[2299] = cin[2237];
assign cj_6144[2300] = cin[4324];
assign cj_6144[2301] = cin[1227];
assign cj_6144[2302] = cin[5234];
assign cj_6144[2303] = cin[4057];
assign cj_6144[2304] = cin[3840];
assign cj_6144[2305] = cin[4583];
assign cj_6144[2306] = cin[142];
assign cj_6144[2307] = cin[2805];
assign cj_6144[2308] = cin[284];
assign cj_6144[2309] = cin[4867];
assign cj_6144[2310] = cin[4266];
assign cj_6144[2311] = cin[4625];
assign cj_6144[2312] = cin[5944];
assign cj_6144[2313] = cin[2079];
assign cj_6144[2314] = cin[5318];
assign cj_6144[2315] = cin[3373];
assign cj_6144[2316] = cin[2388];
assign cj_6144[2317] = cin[2363];
assign cj_6144[2318] = cin[3298];
assign cj_6144[2319] = cin[5193];
assign cj_6144[2320] = cin[1904];
assign cj_6144[2321] = cin[5719];
assign cj_6144[2322] = cin[4350];
assign cj_6144[2323] = cin[3941];
assign cj_6144[2324] = cin[4492];
assign cj_6144[2325] = cin[6003];
assign cj_6144[2326] = cin[2330];
assign cj_6144[2327] = cin[5761];
assign cj_6144[2328] = cin[4008];
assign cj_6144[2329] = cin[3215];
assign cj_6144[2330] = cin[3382];
assign cj_6144[2331] = cin[4509];
assign cj_6144[2332] = cin[452];
assign cj_6144[2333] = cin[3499];
assign cj_6144[2334] = cin[1362];
assign cj_6144[2335] = cin[185];
assign cj_6144[2336] = cin[6112];
assign cj_6144[2337] = cin[711];
assign cj_6144[2338] = cin[2414];
assign cj_6144[2339] = cin[5077];
assign cj_6144[2340] = cin[2556];
assign cj_6144[2341] = cin[995];
assign cj_6144[2342] = cin[394];
assign cj_6144[2343] = cin[753];
assign cj_6144[2344] = cin[2072];
assign cj_6144[2345] = cin[4351];
assign cj_6144[2346] = cin[1446];
assign cj_6144[2347] = cin[5645];
assign cj_6144[2348] = cin[4660];
assign cj_6144[2349] = cin[4635];
assign cj_6144[2350] = cin[5570];
assign cj_6144[2351] = cin[1321];
assign cj_6144[2352] = cin[4176];
assign cj_6144[2353] = cin[1847];
assign cj_6144[2354] = cin[478];
assign cj_6144[2355] = cin[69];
assign cj_6144[2356] = cin[620];
assign cj_6144[2357] = cin[2131];
assign cj_6144[2358] = cin[4602];
assign cj_6144[2359] = cin[1889];
assign cj_6144[2360] = cin[136];
assign cj_6144[2361] = cin[5487];
assign cj_6144[2362] = cin[5654];
assign cj_6144[2363] = cin[637];
assign cj_6144[2364] = cin[2724];
assign cj_6144[2365] = cin[5771];
assign cj_6144[2366] = cin[3634];
assign cj_6144[2367] = cin[2457];
assign cj_6144[2368] = cin[2240];
assign cj_6144[2369] = cin[2983];
assign cj_6144[2370] = cin[4686];
assign cj_6144[2371] = cin[1205];
assign cj_6144[2372] = cin[4828];
assign cj_6144[2373] = cin[3267];
assign cj_6144[2374] = cin[2666];
assign cj_6144[2375] = cin[3025];
assign cj_6144[2376] = cin[4344];
assign cj_6144[2377] = cin[479];
assign cj_6144[2378] = cin[3718];
assign cj_6144[2379] = cin[1773];
assign cj_6144[2380] = cin[788];
assign cj_6144[2381] = cin[763];
assign cj_6144[2382] = cin[1698];
assign cj_6144[2383] = cin[3593];
assign cj_6144[2384] = cin[304];
assign cj_6144[2385] = cin[4119];
assign cj_6144[2386] = cin[2750];
assign cj_6144[2387] = cin[2341];
assign cj_6144[2388] = cin[2892];
assign cj_6144[2389] = cin[4403];
assign cj_6144[2390] = cin[730];
assign cj_6144[2391] = cin[4161];
assign cj_6144[2392] = cin[2408];
assign cj_6144[2393] = cin[1615];
assign cj_6144[2394] = cin[1782];
assign cj_6144[2395] = cin[2909];
assign cj_6144[2396] = cin[4996];
assign cj_6144[2397] = cin[1899];
assign cj_6144[2398] = cin[5906];
assign cj_6144[2399] = cin[4729];
assign cj_6144[2400] = cin[4512];
assign cj_6144[2401] = cin[5255];
assign cj_6144[2402] = cin[814];
assign cj_6144[2403] = cin[3477];
assign cj_6144[2404] = cin[956];
assign cj_6144[2405] = cin[5539];
assign cj_6144[2406] = cin[4938];
assign cj_6144[2407] = cin[5297];
assign cj_6144[2408] = cin[472];
assign cj_6144[2409] = cin[2751];
assign cj_6144[2410] = cin[5990];
assign cj_6144[2411] = cin[4045];
assign cj_6144[2412] = cin[3060];
assign cj_6144[2413] = cin[3035];
assign cj_6144[2414] = cin[3970];
assign cj_6144[2415] = cin[5865];
assign cj_6144[2416] = cin[2576];
assign cj_6144[2417] = cin[247];
assign cj_6144[2418] = cin[5022];
assign cj_6144[2419] = cin[4613];
assign cj_6144[2420] = cin[5164];
assign cj_6144[2421] = cin[531];
assign cj_6144[2422] = cin[3002];
assign cj_6144[2423] = cin[289];
assign cj_6144[2424] = cin[4680];
assign cj_6144[2425] = cin[3887];
assign cj_6144[2426] = cin[4054];
assign cj_6144[2427] = cin[5181];
assign cj_6144[2428] = cin[1124];
assign cj_6144[2429] = cin[4171];
assign cj_6144[2430] = cin[2034];
assign cj_6144[2431] = cin[857];
assign cj_6144[2432] = cin[640];
assign cj_6144[2433] = cin[1383];
assign cj_6144[2434] = cin[3086];
assign cj_6144[2435] = cin[5749];
assign cj_6144[2436] = cin[3228];
assign cj_6144[2437] = cin[1667];
assign cj_6144[2438] = cin[1066];
assign cj_6144[2439] = cin[1425];
assign cj_6144[2440] = cin[2744];
assign cj_6144[2441] = cin[5023];
assign cj_6144[2442] = cin[2118];
assign cj_6144[2443] = cin[173];
assign cj_6144[2444] = cin[5332];
assign cj_6144[2445] = cin[5307];
assign cj_6144[2446] = cin[98];
assign cj_6144[2447] = cin[1993];
assign cj_6144[2448] = cin[4848];
assign cj_6144[2449] = cin[2519];
assign cj_6144[2450] = cin[1150];
assign cj_6144[2451] = cin[741];
assign cj_6144[2452] = cin[1292];
assign cj_6144[2453] = cin[2803];
assign cj_6144[2454] = cin[5274];
assign cj_6144[2455] = cin[2561];
assign cj_6144[2456] = cin[808];
assign cj_6144[2457] = cin[15];
assign cj_6144[2458] = cin[182];
assign cj_6144[2459] = cin[1309];
assign cj_6144[2460] = cin[3396];
assign cj_6144[2461] = cin[299];
assign cj_6144[2462] = cin[4306];
assign cj_6144[2463] = cin[3129];
assign cj_6144[2464] = cin[2912];
assign cj_6144[2465] = cin[3655];
assign cj_6144[2466] = cin[5358];
assign cj_6144[2467] = cin[1877];
assign cj_6144[2468] = cin[5500];
assign cj_6144[2469] = cin[3939];
assign cj_6144[2470] = cin[3338];
assign cj_6144[2471] = cin[3697];
assign cj_6144[2472] = cin[5016];
assign cj_6144[2473] = cin[1151];
assign cj_6144[2474] = cin[4390];
assign cj_6144[2475] = cin[2445];
assign cj_6144[2476] = cin[1460];
assign cj_6144[2477] = cin[1435];
assign cj_6144[2478] = cin[2370];
assign cj_6144[2479] = cin[4265];
assign cj_6144[2480] = cin[976];
assign cj_6144[2481] = cin[4791];
assign cj_6144[2482] = cin[3422];
assign cj_6144[2483] = cin[3013];
assign cj_6144[2484] = cin[3564];
assign cj_6144[2485] = cin[5075];
assign cj_6144[2486] = cin[1402];
assign cj_6144[2487] = cin[4833];
assign cj_6144[2488] = cin[3080];
assign cj_6144[2489] = cin[2287];
assign cj_6144[2490] = cin[2454];
assign cj_6144[2491] = cin[3581];
assign cj_6144[2492] = cin[5668];
assign cj_6144[2493] = cin[2571];
assign cj_6144[2494] = cin[434];
assign cj_6144[2495] = cin[5401];
assign cj_6144[2496] = cin[5184];
assign cj_6144[2497] = cin[5927];
assign cj_6144[2498] = cin[1486];
assign cj_6144[2499] = cin[4149];
assign cj_6144[2500] = cin[1628];
assign cj_6144[2501] = cin[67];
assign cj_6144[2502] = cin[5610];
assign cj_6144[2503] = cin[5969];
assign cj_6144[2504] = cin[1144];
assign cj_6144[2505] = cin[3423];
assign cj_6144[2506] = cin[518];
assign cj_6144[2507] = cin[4717];
assign cj_6144[2508] = cin[3732];
assign cj_6144[2509] = cin[3707];
assign cj_6144[2510] = cin[4642];
assign cj_6144[2511] = cin[393];
assign cj_6144[2512] = cin[3248];
assign cj_6144[2513] = cin[919];
assign cj_6144[2514] = cin[5694];
assign cj_6144[2515] = cin[5285];
assign cj_6144[2516] = cin[5836];
assign cj_6144[2517] = cin[1203];
assign cj_6144[2518] = cin[3674];
assign cj_6144[2519] = cin[961];
assign cj_6144[2520] = cin[5352];
assign cj_6144[2521] = cin[4559];
assign cj_6144[2522] = cin[4726];
assign cj_6144[2523] = cin[5853];
assign cj_6144[2524] = cin[1796];
assign cj_6144[2525] = cin[4843];
assign cj_6144[2526] = cin[2706];
assign cj_6144[2527] = cin[1529];
assign cj_6144[2528] = cin[1312];
assign cj_6144[2529] = cin[2055];
assign cj_6144[2530] = cin[3758];
assign cj_6144[2531] = cin[277];
assign cj_6144[2532] = cin[3900];
assign cj_6144[2533] = cin[2339];
assign cj_6144[2534] = cin[1738];
assign cj_6144[2535] = cin[2097];
assign cj_6144[2536] = cin[3416];
assign cj_6144[2537] = cin[5695];
assign cj_6144[2538] = cin[2790];
assign cj_6144[2539] = cin[845];
assign cj_6144[2540] = cin[6004];
assign cj_6144[2541] = cin[5979];
assign cj_6144[2542] = cin[770];
assign cj_6144[2543] = cin[2665];
assign cj_6144[2544] = cin[5520];
assign cj_6144[2545] = cin[3191];
assign cj_6144[2546] = cin[1822];
assign cj_6144[2547] = cin[1413];
assign cj_6144[2548] = cin[1964];
assign cj_6144[2549] = cin[3475];
assign cj_6144[2550] = cin[5946];
assign cj_6144[2551] = cin[3233];
assign cj_6144[2552] = cin[1480];
assign cj_6144[2553] = cin[687];
assign cj_6144[2554] = cin[854];
assign cj_6144[2555] = cin[1981];
assign cj_6144[2556] = cin[4068];
assign cj_6144[2557] = cin[971];
assign cj_6144[2558] = cin[4978];
assign cj_6144[2559] = cin[3801];
assign cj_6144[2560] = cin[3584];
assign cj_6144[2561] = cin[4327];
assign cj_6144[2562] = cin[6030];
assign cj_6144[2563] = cin[2549];
assign cj_6144[2564] = cin[28];
assign cj_6144[2565] = cin[4611];
assign cj_6144[2566] = cin[4010];
assign cj_6144[2567] = cin[4369];
assign cj_6144[2568] = cin[5688];
assign cj_6144[2569] = cin[1823];
assign cj_6144[2570] = cin[5062];
assign cj_6144[2571] = cin[3117];
assign cj_6144[2572] = cin[2132];
assign cj_6144[2573] = cin[2107];
assign cj_6144[2574] = cin[3042];
assign cj_6144[2575] = cin[4937];
assign cj_6144[2576] = cin[1648];
assign cj_6144[2577] = cin[5463];
assign cj_6144[2578] = cin[4094];
assign cj_6144[2579] = cin[3685];
assign cj_6144[2580] = cin[4236];
assign cj_6144[2581] = cin[5747];
assign cj_6144[2582] = cin[2074];
assign cj_6144[2583] = cin[5505];
assign cj_6144[2584] = cin[3752];
assign cj_6144[2585] = cin[2959];
assign cj_6144[2586] = cin[3126];
assign cj_6144[2587] = cin[4253];
assign cj_6144[2588] = cin[196];
assign cj_6144[2589] = cin[3243];
assign cj_6144[2590] = cin[1106];
assign cj_6144[2591] = cin[6073];
assign cj_6144[2592] = cin[5856];
assign cj_6144[2593] = cin[455];
assign cj_6144[2594] = cin[2158];
assign cj_6144[2595] = cin[4821];
assign cj_6144[2596] = cin[2300];
assign cj_6144[2597] = cin[739];
assign cj_6144[2598] = cin[138];
assign cj_6144[2599] = cin[497];
assign cj_6144[2600] = cin[1816];
assign cj_6144[2601] = cin[4095];
assign cj_6144[2602] = cin[1190];
assign cj_6144[2603] = cin[5389];
assign cj_6144[2604] = cin[4404];
assign cj_6144[2605] = cin[4379];
assign cj_6144[2606] = cin[5314];
assign cj_6144[2607] = cin[1065];
assign cj_6144[2608] = cin[3920];
assign cj_6144[2609] = cin[1591];
assign cj_6144[2610] = cin[222];
assign cj_6144[2611] = cin[5957];
assign cj_6144[2612] = cin[364];
assign cj_6144[2613] = cin[1875];
assign cj_6144[2614] = cin[4346];
assign cj_6144[2615] = cin[1633];
assign cj_6144[2616] = cin[6024];
assign cj_6144[2617] = cin[5231];
assign cj_6144[2618] = cin[5398];
assign cj_6144[2619] = cin[381];
assign cj_6144[2620] = cin[2468];
assign cj_6144[2621] = cin[5515];
assign cj_6144[2622] = cin[3378];
assign cj_6144[2623] = cin[2201];
assign cj_6144[2624] = cin[1984];
assign cj_6144[2625] = cin[2727];
assign cj_6144[2626] = cin[4430];
assign cj_6144[2627] = cin[949];
assign cj_6144[2628] = cin[4572];
assign cj_6144[2629] = cin[3011];
assign cj_6144[2630] = cin[2410];
assign cj_6144[2631] = cin[2769];
assign cj_6144[2632] = cin[4088];
assign cj_6144[2633] = cin[223];
assign cj_6144[2634] = cin[3462];
assign cj_6144[2635] = cin[1517];
assign cj_6144[2636] = cin[532];
assign cj_6144[2637] = cin[507];
assign cj_6144[2638] = cin[1442];
assign cj_6144[2639] = cin[3337];
assign cj_6144[2640] = cin[48];
assign cj_6144[2641] = cin[3863];
assign cj_6144[2642] = cin[2494];
assign cj_6144[2643] = cin[2085];
assign cj_6144[2644] = cin[2636];
assign cj_6144[2645] = cin[4147];
assign cj_6144[2646] = cin[474];
assign cj_6144[2647] = cin[3905];
assign cj_6144[2648] = cin[2152];
assign cj_6144[2649] = cin[1359];
assign cj_6144[2650] = cin[1526];
assign cj_6144[2651] = cin[2653];
assign cj_6144[2652] = cin[4740];
assign cj_6144[2653] = cin[1643];
assign cj_6144[2654] = cin[5650];
assign cj_6144[2655] = cin[4473];
assign cj_6144[2656] = cin[4256];
assign cj_6144[2657] = cin[4999];
assign cj_6144[2658] = cin[558];
assign cj_6144[2659] = cin[3221];
assign cj_6144[2660] = cin[700];
assign cj_6144[2661] = cin[5283];
assign cj_6144[2662] = cin[4682];
assign cj_6144[2663] = cin[5041];
assign cj_6144[2664] = cin[216];
assign cj_6144[2665] = cin[2495];
assign cj_6144[2666] = cin[5734];
assign cj_6144[2667] = cin[3789];
assign cj_6144[2668] = cin[2804];
assign cj_6144[2669] = cin[2779];
assign cj_6144[2670] = cin[3714];
assign cj_6144[2671] = cin[5609];
assign cj_6144[2672] = cin[2320];
assign cj_6144[2673] = cin[6135];
assign cj_6144[2674] = cin[4766];
assign cj_6144[2675] = cin[4357];
assign cj_6144[2676] = cin[4908];
assign cj_6144[2677] = cin[275];
assign cj_6144[2678] = cin[2746];
assign cj_6144[2679] = cin[33];
assign cj_6144[2680] = cin[4424];
assign cj_6144[2681] = cin[3631];
assign cj_6144[2682] = cin[3798];
assign cj_6144[2683] = cin[4925];
assign cj_6144[2684] = cin[868];
assign cj_6144[2685] = cin[3915];
assign cj_6144[2686] = cin[1778];
assign cj_6144[2687] = cin[601];
assign cj_6144[2688] = cin[384];
assign cj_6144[2689] = cin[1127];
assign cj_6144[2690] = cin[2830];
assign cj_6144[2691] = cin[5493];
assign cj_6144[2692] = cin[2972];
assign cj_6144[2693] = cin[1411];
assign cj_6144[2694] = cin[810];
assign cj_6144[2695] = cin[1169];
assign cj_6144[2696] = cin[2488];
assign cj_6144[2697] = cin[4767];
assign cj_6144[2698] = cin[1862];
assign cj_6144[2699] = cin[6061];
assign cj_6144[2700] = cin[5076];
assign cj_6144[2701] = cin[5051];
assign cj_6144[2702] = cin[5986];
assign cj_6144[2703] = cin[1737];
assign cj_6144[2704] = cin[4592];
assign cj_6144[2705] = cin[2263];
assign cj_6144[2706] = cin[894];
assign cj_6144[2707] = cin[485];
assign cj_6144[2708] = cin[1036];
assign cj_6144[2709] = cin[2547];
assign cj_6144[2710] = cin[5018];
assign cj_6144[2711] = cin[2305];
assign cj_6144[2712] = cin[552];
assign cj_6144[2713] = cin[5903];
assign cj_6144[2714] = cin[6070];
assign cj_6144[2715] = cin[1053];
assign cj_6144[2716] = cin[3140];
assign cj_6144[2717] = cin[43];
assign cj_6144[2718] = cin[4050];
assign cj_6144[2719] = cin[2873];
assign cj_6144[2720] = cin[2656];
assign cj_6144[2721] = cin[3399];
assign cj_6144[2722] = cin[5102];
assign cj_6144[2723] = cin[1621];
assign cj_6144[2724] = cin[5244];
assign cj_6144[2725] = cin[3683];
assign cj_6144[2726] = cin[3082];
assign cj_6144[2727] = cin[3441];
assign cj_6144[2728] = cin[4760];
assign cj_6144[2729] = cin[895];
assign cj_6144[2730] = cin[4134];
assign cj_6144[2731] = cin[2189];
assign cj_6144[2732] = cin[1204];
assign cj_6144[2733] = cin[1179];
assign cj_6144[2734] = cin[2114];
assign cj_6144[2735] = cin[4009];
assign cj_6144[2736] = cin[720];
assign cj_6144[2737] = cin[4535];
assign cj_6144[2738] = cin[3166];
assign cj_6144[2739] = cin[2757];
assign cj_6144[2740] = cin[3308];
assign cj_6144[2741] = cin[4819];
assign cj_6144[2742] = cin[1146];
assign cj_6144[2743] = cin[4577];
assign cj_6144[2744] = cin[2824];
assign cj_6144[2745] = cin[2031];
assign cj_6144[2746] = cin[2198];
assign cj_6144[2747] = cin[3325];
assign cj_6144[2748] = cin[5412];
assign cj_6144[2749] = cin[2315];
assign cj_6144[2750] = cin[178];
assign cj_6144[2751] = cin[5145];
assign cj_6144[2752] = cin[4928];
assign cj_6144[2753] = cin[5671];
assign cj_6144[2754] = cin[1230];
assign cj_6144[2755] = cin[3893];
assign cj_6144[2756] = cin[1372];
assign cj_6144[2757] = cin[5955];
assign cj_6144[2758] = cin[5354];
assign cj_6144[2759] = cin[5713];
assign cj_6144[2760] = cin[888];
assign cj_6144[2761] = cin[3167];
assign cj_6144[2762] = cin[262];
assign cj_6144[2763] = cin[4461];
assign cj_6144[2764] = cin[3476];
assign cj_6144[2765] = cin[3451];
assign cj_6144[2766] = cin[4386];
assign cj_6144[2767] = cin[137];
assign cj_6144[2768] = cin[2992];
assign cj_6144[2769] = cin[663];
assign cj_6144[2770] = cin[5438];
assign cj_6144[2771] = cin[5029];
assign cj_6144[2772] = cin[5580];
assign cj_6144[2773] = cin[947];
assign cj_6144[2774] = cin[3418];
assign cj_6144[2775] = cin[705];
assign cj_6144[2776] = cin[5096];
assign cj_6144[2777] = cin[4303];
assign cj_6144[2778] = cin[4470];
assign cj_6144[2779] = cin[5597];
assign cj_6144[2780] = cin[1540];
assign cj_6144[2781] = cin[4587];
assign cj_6144[2782] = cin[2450];
assign cj_6144[2783] = cin[1273];
assign cj_6144[2784] = cin[1056];
assign cj_6144[2785] = cin[1799];
assign cj_6144[2786] = cin[3502];
assign cj_6144[2787] = cin[21];
assign cj_6144[2788] = cin[3644];
assign cj_6144[2789] = cin[2083];
assign cj_6144[2790] = cin[1482];
assign cj_6144[2791] = cin[1841];
assign cj_6144[2792] = cin[3160];
assign cj_6144[2793] = cin[5439];
assign cj_6144[2794] = cin[2534];
assign cj_6144[2795] = cin[589];
assign cj_6144[2796] = cin[5748];
assign cj_6144[2797] = cin[5723];
assign cj_6144[2798] = cin[514];
assign cj_6144[2799] = cin[2409];
assign cj_6144[2800] = cin[5264];
assign cj_6144[2801] = cin[2935];
assign cj_6144[2802] = cin[1566];
assign cj_6144[2803] = cin[1157];
assign cj_6144[2804] = cin[1708];
assign cj_6144[2805] = cin[3219];
assign cj_6144[2806] = cin[5690];
assign cj_6144[2807] = cin[2977];
assign cj_6144[2808] = cin[1224];
assign cj_6144[2809] = cin[431];
assign cj_6144[2810] = cin[598];
assign cj_6144[2811] = cin[1725];
assign cj_6144[2812] = cin[3812];
assign cj_6144[2813] = cin[715];
assign cj_6144[2814] = cin[4722];
assign cj_6144[2815] = cin[3545];
assign cj_6144[2816] = cin[3328];
assign cj_6144[2817] = cin[4071];
assign cj_6144[2818] = cin[5774];
assign cj_6144[2819] = cin[2293];
assign cj_6144[2820] = cin[5916];
assign cj_6144[2821] = cin[4355];
assign cj_6144[2822] = cin[3754];
assign cj_6144[2823] = cin[4113];
assign cj_6144[2824] = cin[5432];
assign cj_6144[2825] = cin[1567];
assign cj_6144[2826] = cin[4806];
assign cj_6144[2827] = cin[2861];
assign cj_6144[2828] = cin[1876];
assign cj_6144[2829] = cin[1851];
assign cj_6144[2830] = cin[2786];
assign cj_6144[2831] = cin[4681];
assign cj_6144[2832] = cin[1392];
assign cj_6144[2833] = cin[5207];
assign cj_6144[2834] = cin[3838];
assign cj_6144[2835] = cin[3429];
assign cj_6144[2836] = cin[3980];
assign cj_6144[2837] = cin[5491];
assign cj_6144[2838] = cin[1818];
assign cj_6144[2839] = cin[5249];
assign cj_6144[2840] = cin[3496];
assign cj_6144[2841] = cin[2703];
assign cj_6144[2842] = cin[2870];
assign cj_6144[2843] = cin[3997];
assign cj_6144[2844] = cin[6084];
assign cj_6144[2845] = cin[2987];
assign cj_6144[2846] = cin[850];
assign cj_6144[2847] = cin[5817];
assign cj_6144[2848] = cin[5600];
assign cj_6144[2849] = cin[199];
assign cj_6144[2850] = cin[1902];
assign cj_6144[2851] = cin[4565];
assign cj_6144[2852] = cin[2044];
assign cj_6144[2853] = cin[483];
assign cj_6144[2854] = cin[6026];
assign cj_6144[2855] = cin[241];
assign cj_6144[2856] = cin[1560];
assign cj_6144[2857] = cin[3839];
assign cj_6144[2858] = cin[934];
assign cj_6144[2859] = cin[5133];
assign cj_6144[2860] = cin[4148];
assign cj_6144[2861] = cin[4123];
assign cj_6144[2862] = cin[5058];
assign cj_6144[2863] = cin[809];
assign cj_6144[2864] = cin[3664];
assign cj_6144[2865] = cin[1335];
assign cj_6144[2866] = cin[6110];
assign cj_6144[2867] = cin[5701];
assign cj_6144[2868] = cin[108];
assign cj_6144[2869] = cin[1619];
assign cj_6144[2870] = cin[4090];
assign cj_6144[2871] = cin[1377];
assign cj_6144[2872] = cin[5768];
assign cj_6144[2873] = cin[4975];
assign cj_6144[2874] = cin[5142];
assign cj_6144[2875] = cin[125];
assign cj_6144[2876] = cin[2212];
assign cj_6144[2877] = cin[5259];
assign cj_6144[2878] = cin[3122];
assign cj_6144[2879] = cin[1945];
assign cj_6144[2880] = cin[1728];
assign cj_6144[2881] = cin[2471];
assign cj_6144[2882] = cin[4174];
assign cj_6144[2883] = cin[693];
assign cj_6144[2884] = cin[4316];
assign cj_6144[2885] = cin[2755];
assign cj_6144[2886] = cin[2154];
assign cj_6144[2887] = cin[2513];
assign cj_6144[2888] = cin[3832];
assign cj_6144[2889] = cin[6111];
assign cj_6144[2890] = cin[3206];
assign cj_6144[2891] = cin[1261];
assign cj_6144[2892] = cin[276];
assign cj_6144[2893] = cin[251];
assign cj_6144[2894] = cin[1186];
assign cj_6144[2895] = cin[3081];
assign cj_6144[2896] = cin[5936];
assign cj_6144[2897] = cin[3607];
assign cj_6144[2898] = cin[2238];
assign cj_6144[2899] = cin[1829];
assign cj_6144[2900] = cin[2380];
assign cj_6144[2901] = cin[3891];
assign cj_6144[2902] = cin[218];
assign cj_6144[2903] = cin[3649];
assign cj_6144[2904] = cin[1896];
assign cj_6144[2905] = cin[1103];
assign cj_6144[2906] = cin[1270];
assign cj_6144[2907] = cin[2397];
assign cj_6144[2908] = cin[4484];
assign cj_6144[2909] = cin[1387];
assign cj_6144[2910] = cin[5394];
assign cj_6144[2911] = cin[4217];
assign cj_6144[2912] = cin[4000];
assign cj_6144[2913] = cin[4743];
assign cj_6144[2914] = cin[302];
assign cj_6144[2915] = cin[2965];
assign cj_6144[2916] = cin[444];
assign cj_6144[2917] = cin[5027];
assign cj_6144[2918] = cin[4426];
assign cj_6144[2919] = cin[4785];
assign cj_6144[2920] = cin[6104];
assign cj_6144[2921] = cin[2239];
assign cj_6144[2922] = cin[5478];
assign cj_6144[2923] = cin[3533];
assign cj_6144[2924] = cin[2548];
assign cj_6144[2925] = cin[2523];
assign cj_6144[2926] = cin[3458];
assign cj_6144[2927] = cin[5353];
assign cj_6144[2928] = cin[2064];
assign cj_6144[2929] = cin[5879];
assign cj_6144[2930] = cin[4510];
assign cj_6144[2931] = cin[4101];
assign cj_6144[2932] = cin[4652];
assign cj_6144[2933] = cin[19];
assign cj_6144[2934] = cin[2490];
assign cj_6144[2935] = cin[5921];
assign cj_6144[2936] = cin[4168];
assign cj_6144[2937] = cin[3375];
assign cj_6144[2938] = cin[3542];
assign cj_6144[2939] = cin[4669];
assign cj_6144[2940] = cin[612];
assign cj_6144[2941] = cin[3659];
assign cj_6144[2942] = cin[1522];
assign cj_6144[2943] = cin[345];
assign cj_6144[2944] = cin[128];
assign cj_6144[2945] = cin[871];
assign cj_6144[2946] = cin[2574];
assign cj_6144[2947] = cin[5237];
assign cj_6144[2948] = cin[2716];
assign cj_6144[2949] = cin[1155];
assign cj_6144[2950] = cin[554];
assign cj_6144[2951] = cin[913];
assign cj_6144[2952] = cin[2232];
assign cj_6144[2953] = cin[4511];
assign cj_6144[2954] = cin[1606];
assign cj_6144[2955] = cin[5805];
assign cj_6144[2956] = cin[4820];
assign cj_6144[2957] = cin[4795];
assign cj_6144[2958] = cin[5730];
assign cj_6144[2959] = cin[1481];
assign cj_6144[2960] = cin[4336];
assign cj_6144[2961] = cin[2007];
assign cj_6144[2962] = cin[638];
assign cj_6144[2963] = cin[229];
assign cj_6144[2964] = cin[780];
assign cj_6144[2965] = cin[2291];
assign cj_6144[2966] = cin[4762];
assign cj_6144[2967] = cin[2049];
assign cj_6144[2968] = cin[296];
assign cj_6144[2969] = cin[5647];
assign cj_6144[2970] = cin[5814];
assign cj_6144[2971] = cin[797];
assign cj_6144[2972] = cin[2884];
assign cj_6144[2973] = cin[5931];
assign cj_6144[2974] = cin[3794];
assign cj_6144[2975] = cin[2617];
assign cj_6144[2976] = cin[2400];
assign cj_6144[2977] = cin[3143];
assign cj_6144[2978] = cin[4846];
assign cj_6144[2979] = cin[1365];
assign cj_6144[2980] = cin[4988];
assign cj_6144[2981] = cin[3427];
assign cj_6144[2982] = cin[2826];
assign cj_6144[2983] = cin[3185];
assign cj_6144[2984] = cin[4504];
assign cj_6144[2985] = cin[639];
assign cj_6144[2986] = cin[3878];
assign cj_6144[2987] = cin[1933];
assign cj_6144[2988] = cin[948];
assign cj_6144[2989] = cin[923];
assign cj_6144[2990] = cin[1858];
assign cj_6144[2991] = cin[3753];
assign cj_6144[2992] = cin[464];
assign cj_6144[2993] = cin[4279];
assign cj_6144[2994] = cin[2910];
assign cj_6144[2995] = cin[2501];
assign cj_6144[2996] = cin[3052];
assign cj_6144[2997] = cin[4563];
assign cj_6144[2998] = cin[890];
assign cj_6144[2999] = cin[4321];
assign cj_6144[3000] = cin[2568];
assign cj_6144[3001] = cin[1775];
assign cj_6144[3002] = cin[1942];
assign cj_6144[3003] = cin[3069];
assign cj_6144[3004] = cin[5156];
assign cj_6144[3005] = cin[2059];
assign cj_6144[3006] = cin[6066];
assign cj_6144[3007] = cin[4889];
assign cj_6144[3008] = cin[4672];
assign cj_6144[3009] = cin[5415];
assign cj_6144[3010] = cin[974];
assign cj_6144[3011] = cin[3637];
assign cj_6144[3012] = cin[1116];
assign cj_6144[3013] = cin[5699];
assign cj_6144[3014] = cin[5098];
assign cj_6144[3015] = cin[5457];
assign cj_6144[3016] = cin[632];
assign cj_6144[3017] = cin[2911];
assign cj_6144[3018] = cin[6];
assign cj_6144[3019] = cin[4205];
assign cj_6144[3020] = cin[3220];
assign cj_6144[3021] = cin[3195];
assign cj_6144[3022] = cin[4130];
assign cj_6144[3023] = cin[6025];
assign cj_6144[3024] = cin[2736];
assign cj_6144[3025] = cin[407];
assign cj_6144[3026] = cin[5182];
assign cj_6144[3027] = cin[4773];
assign cj_6144[3028] = cin[5324];
assign cj_6144[3029] = cin[691];
assign cj_6144[3030] = cin[3162];
assign cj_6144[3031] = cin[449];
assign cj_6144[3032] = cin[4840];
assign cj_6144[3033] = cin[4047];
assign cj_6144[3034] = cin[4214];
assign cj_6144[3035] = cin[5341];
assign cj_6144[3036] = cin[1284];
assign cj_6144[3037] = cin[4331];
assign cj_6144[3038] = cin[2194];
assign cj_6144[3039] = cin[1017];
assign cj_6144[3040] = cin[800];
assign cj_6144[3041] = cin[1543];
assign cj_6144[3042] = cin[3246];
assign cj_6144[3043] = cin[5909];
assign cj_6144[3044] = cin[3388];
assign cj_6144[3045] = cin[1827];
assign cj_6144[3046] = cin[1226];
assign cj_6144[3047] = cin[1585];
assign cj_6144[3048] = cin[2904];
assign cj_6144[3049] = cin[5183];
assign cj_6144[3050] = cin[2278];
assign cj_6144[3051] = cin[333];
assign cj_6144[3052] = cin[5492];
assign cj_6144[3053] = cin[5467];
assign cj_6144[3054] = cin[258];
assign cj_6144[3055] = cin[2153];
assign cj_6144[3056] = cin[5008];
assign cj_6144[3057] = cin[2679];
assign cj_6144[3058] = cin[1310];
assign cj_6144[3059] = cin[901];
assign cj_6144[3060] = cin[1452];
assign cj_6144[3061] = cin[2963];
assign cj_6144[3062] = cin[5434];
assign cj_6144[3063] = cin[2721];
assign cj_6144[3064] = cin[968];
assign cj_6144[3065] = cin[175];
assign cj_6144[3066] = cin[342];
assign cj_6144[3067] = cin[1469];
assign cj_6144[3068] = cin[3556];
assign cj_6144[3069] = cin[459];
assign cj_6144[3070] = cin[4466];
assign cj_6144[3071] = cin[3289];
assign cj_6144[3072] = cin[3072];
assign cj_6144[3073] = cin[3815];
assign cj_6144[3074] = cin[5518];
assign cj_6144[3075] = cin[2037];
assign cj_6144[3076] = cin[5660];
assign cj_6144[3077] = cin[4099];
assign cj_6144[3078] = cin[3498];
assign cj_6144[3079] = cin[3857];
assign cj_6144[3080] = cin[5176];
assign cj_6144[3081] = cin[1311];
assign cj_6144[3082] = cin[4550];
assign cj_6144[3083] = cin[2605];
assign cj_6144[3084] = cin[1620];
assign cj_6144[3085] = cin[1595];
assign cj_6144[3086] = cin[2530];
assign cj_6144[3087] = cin[4425];
assign cj_6144[3088] = cin[1136];
assign cj_6144[3089] = cin[4951];
assign cj_6144[3090] = cin[3582];
assign cj_6144[3091] = cin[3173];
assign cj_6144[3092] = cin[3724];
assign cj_6144[3093] = cin[5235];
assign cj_6144[3094] = cin[1562];
assign cj_6144[3095] = cin[4993];
assign cj_6144[3096] = cin[3240];
assign cj_6144[3097] = cin[2447];
assign cj_6144[3098] = cin[2614];
assign cj_6144[3099] = cin[3741];
assign cj_6144[3100] = cin[5828];
assign cj_6144[3101] = cin[2731];
assign cj_6144[3102] = cin[594];
assign cj_6144[3103] = cin[5561];
assign cj_6144[3104] = cin[5344];
assign cj_6144[3105] = cin[6087];
assign cj_6144[3106] = cin[1646];
assign cj_6144[3107] = cin[4309];
assign cj_6144[3108] = cin[1788];
assign cj_6144[3109] = cin[227];
assign cj_6144[3110] = cin[5770];
assign cj_6144[3111] = cin[6129];
assign cj_6144[3112] = cin[1304];
assign cj_6144[3113] = cin[3583];
assign cj_6144[3114] = cin[678];
assign cj_6144[3115] = cin[4877];
assign cj_6144[3116] = cin[3892];
assign cj_6144[3117] = cin[3867];
assign cj_6144[3118] = cin[4802];
assign cj_6144[3119] = cin[553];
assign cj_6144[3120] = cin[3408];
assign cj_6144[3121] = cin[1079];
assign cj_6144[3122] = cin[5854];
assign cj_6144[3123] = cin[5445];
assign cj_6144[3124] = cin[5996];
assign cj_6144[3125] = cin[1363];
assign cj_6144[3126] = cin[3834];
assign cj_6144[3127] = cin[1121];
assign cj_6144[3128] = cin[5512];
assign cj_6144[3129] = cin[4719];
assign cj_6144[3130] = cin[4886];
assign cj_6144[3131] = cin[6013];
assign cj_6144[3132] = cin[1956];
assign cj_6144[3133] = cin[5003];
assign cj_6144[3134] = cin[2866];
assign cj_6144[3135] = cin[1689];
assign cj_6144[3136] = cin[1472];
assign cj_6144[3137] = cin[2215];
assign cj_6144[3138] = cin[3918];
assign cj_6144[3139] = cin[437];
assign cj_6144[3140] = cin[4060];
assign cj_6144[3141] = cin[2499];
assign cj_6144[3142] = cin[1898];
assign cj_6144[3143] = cin[2257];
assign cj_6144[3144] = cin[3576];
assign cj_6144[3145] = cin[5855];
assign cj_6144[3146] = cin[2950];
assign cj_6144[3147] = cin[1005];
assign cj_6144[3148] = cin[20];
assign cj_6144[3149] = cin[6139];
assign cj_6144[3150] = cin[930];
assign cj_6144[3151] = cin[2825];
assign cj_6144[3152] = cin[5680];
assign cj_6144[3153] = cin[3351];
assign cj_6144[3154] = cin[1982];
assign cj_6144[3155] = cin[1573];
assign cj_6144[3156] = cin[2124];
assign cj_6144[3157] = cin[3635];
assign cj_6144[3158] = cin[6106];
assign cj_6144[3159] = cin[3393];
assign cj_6144[3160] = cin[1640];
assign cj_6144[3161] = cin[847];
assign cj_6144[3162] = cin[1014];
assign cj_6144[3163] = cin[2141];
assign cj_6144[3164] = cin[4228];
assign cj_6144[3165] = cin[1131];
assign cj_6144[3166] = cin[5138];
assign cj_6144[3167] = cin[3961];
assign cj_6144[3168] = cin[3744];
assign cj_6144[3169] = cin[4487];
assign cj_6144[3170] = cin[46];
assign cj_6144[3171] = cin[2709];
assign cj_6144[3172] = cin[188];
assign cj_6144[3173] = cin[4771];
assign cj_6144[3174] = cin[4170];
assign cj_6144[3175] = cin[4529];
assign cj_6144[3176] = cin[5848];
assign cj_6144[3177] = cin[1983];
assign cj_6144[3178] = cin[5222];
assign cj_6144[3179] = cin[3277];
assign cj_6144[3180] = cin[2292];
assign cj_6144[3181] = cin[2267];
assign cj_6144[3182] = cin[3202];
assign cj_6144[3183] = cin[5097];
assign cj_6144[3184] = cin[1808];
assign cj_6144[3185] = cin[5623];
assign cj_6144[3186] = cin[4254];
assign cj_6144[3187] = cin[3845];
assign cj_6144[3188] = cin[4396];
assign cj_6144[3189] = cin[5907];
assign cj_6144[3190] = cin[2234];
assign cj_6144[3191] = cin[5665];
assign cj_6144[3192] = cin[3912];
assign cj_6144[3193] = cin[3119];
assign cj_6144[3194] = cin[3286];
assign cj_6144[3195] = cin[4413];
assign cj_6144[3196] = cin[356];
assign cj_6144[3197] = cin[3403];
assign cj_6144[3198] = cin[1266];
assign cj_6144[3199] = cin[89];
assign cj_6144[3200] = cin[6016];
assign cj_6144[3201] = cin[615];
assign cj_6144[3202] = cin[2318];
assign cj_6144[3203] = cin[4981];
assign cj_6144[3204] = cin[2460];
assign cj_6144[3205] = cin[899];
assign cj_6144[3206] = cin[298];
assign cj_6144[3207] = cin[657];
assign cj_6144[3208] = cin[1976];
assign cj_6144[3209] = cin[4255];
assign cj_6144[3210] = cin[1350];
assign cj_6144[3211] = cin[5549];
assign cj_6144[3212] = cin[4564];
assign cj_6144[3213] = cin[4539];
assign cj_6144[3214] = cin[5474];
assign cj_6144[3215] = cin[1225];
assign cj_6144[3216] = cin[4080];
assign cj_6144[3217] = cin[1751];
assign cj_6144[3218] = cin[382];
assign cj_6144[3219] = cin[6117];
assign cj_6144[3220] = cin[524];
assign cj_6144[3221] = cin[2035];
assign cj_6144[3222] = cin[4506];
assign cj_6144[3223] = cin[1793];
assign cj_6144[3224] = cin[40];
assign cj_6144[3225] = cin[5391];
assign cj_6144[3226] = cin[5558];
assign cj_6144[3227] = cin[541];
assign cj_6144[3228] = cin[2628];
assign cj_6144[3229] = cin[5675];
assign cj_6144[3230] = cin[3538];
assign cj_6144[3231] = cin[2361];
assign cj_6144[3232] = cin[2144];
assign cj_6144[3233] = cin[2887];
assign cj_6144[3234] = cin[4590];
assign cj_6144[3235] = cin[1109];
assign cj_6144[3236] = cin[4732];
assign cj_6144[3237] = cin[3171];
assign cj_6144[3238] = cin[2570];
assign cj_6144[3239] = cin[2929];
assign cj_6144[3240] = cin[4248];
assign cj_6144[3241] = cin[383];
assign cj_6144[3242] = cin[3622];
assign cj_6144[3243] = cin[1677];
assign cj_6144[3244] = cin[692];
assign cj_6144[3245] = cin[667];
assign cj_6144[3246] = cin[1602];
assign cj_6144[3247] = cin[3497];
assign cj_6144[3248] = cin[208];
assign cj_6144[3249] = cin[4023];
assign cj_6144[3250] = cin[2654];
assign cj_6144[3251] = cin[2245];
assign cj_6144[3252] = cin[2796];
assign cj_6144[3253] = cin[4307];
assign cj_6144[3254] = cin[634];
assign cj_6144[3255] = cin[4065];
assign cj_6144[3256] = cin[2312];
assign cj_6144[3257] = cin[1519];
assign cj_6144[3258] = cin[1686];
assign cj_6144[3259] = cin[2813];
assign cj_6144[3260] = cin[4900];
assign cj_6144[3261] = cin[1803];
assign cj_6144[3262] = cin[5810];
assign cj_6144[3263] = cin[4633];
assign cj_6144[3264] = cin[4416];
assign cj_6144[3265] = cin[5159];
assign cj_6144[3266] = cin[718];
assign cj_6144[3267] = cin[3381];
assign cj_6144[3268] = cin[860];
assign cj_6144[3269] = cin[5443];
assign cj_6144[3270] = cin[4842];
assign cj_6144[3271] = cin[5201];
assign cj_6144[3272] = cin[376];
assign cj_6144[3273] = cin[2655];
assign cj_6144[3274] = cin[5894];
assign cj_6144[3275] = cin[3949];
assign cj_6144[3276] = cin[2964];
assign cj_6144[3277] = cin[2939];
assign cj_6144[3278] = cin[3874];
assign cj_6144[3279] = cin[5769];
assign cj_6144[3280] = cin[2480];
assign cj_6144[3281] = cin[151];
assign cj_6144[3282] = cin[4926];
assign cj_6144[3283] = cin[4517];
assign cj_6144[3284] = cin[5068];
assign cj_6144[3285] = cin[435];
assign cj_6144[3286] = cin[2906];
assign cj_6144[3287] = cin[193];
assign cj_6144[3288] = cin[4584];
assign cj_6144[3289] = cin[3791];
assign cj_6144[3290] = cin[3958];
assign cj_6144[3291] = cin[5085];
assign cj_6144[3292] = cin[1028];
assign cj_6144[3293] = cin[4075];
assign cj_6144[3294] = cin[1938];
assign cj_6144[3295] = cin[761];
assign cj_6144[3296] = cin[544];
assign cj_6144[3297] = cin[1287];
assign cj_6144[3298] = cin[2990];
assign cj_6144[3299] = cin[5653];
assign cj_6144[3300] = cin[3132];
assign cj_6144[3301] = cin[1571];
assign cj_6144[3302] = cin[970];
assign cj_6144[3303] = cin[1329];
assign cj_6144[3304] = cin[2648];
assign cj_6144[3305] = cin[4927];
assign cj_6144[3306] = cin[2022];
assign cj_6144[3307] = cin[77];
assign cj_6144[3308] = cin[5236];
assign cj_6144[3309] = cin[5211];
assign cj_6144[3310] = cin[2];
assign cj_6144[3311] = cin[1897];
assign cj_6144[3312] = cin[4752];
assign cj_6144[3313] = cin[2423];
assign cj_6144[3314] = cin[1054];
assign cj_6144[3315] = cin[645];
assign cj_6144[3316] = cin[1196];
assign cj_6144[3317] = cin[2707];
assign cj_6144[3318] = cin[5178];
assign cj_6144[3319] = cin[2465];
assign cj_6144[3320] = cin[712];
assign cj_6144[3321] = cin[6063];
assign cj_6144[3322] = cin[86];
assign cj_6144[3323] = cin[1213];
assign cj_6144[3324] = cin[3300];
assign cj_6144[3325] = cin[203];
assign cj_6144[3326] = cin[4210];
assign cj_6144[3327] = cin[3033];
assign cj_6144[3328] = cin[2816];
assign cj_6144[3329] = cin[3559];
assign cj_6144[3330] = cin[5262];
assign cj_6144[3331] = cin[1781];
assign cj_6144[3332] = cin[5404];
assign cj_6144[3333] = cin[3843];
assign cj_6144[3334] = cin[3242];
assign cj_6144[3335] = cin[3601];
assign cj_6144[3336] = cin[4920];
assign cj_6144[3337] = cin[1055];
assign cj_6144[3338] = cin[4294];
assign cj_6144[3339] = cin[2349];
assign cj_6144[3340] = cin[1364];
assign cj_6144[3341] = cin[1339];
assign cj_6144[3342] = cin[2274];
assign cj_6144[3343] = cin[4169];
assign cj_6144[3344] = cin[880];
assign cj_6144[3345] = cin[4695];
assign cj_6144[3346] = cin[3326];
assign cj_6144[3347] = cin[2917];
assign cj_6144[3348] = cin[3468];
assign cj_6144[3349] = cin[4979];
assign cj_6144[3350] = cin[1306];
assign cj_6144[3351] = cin[4737];
assign cj_6144[3352] = cin[2984];
assign cj_6144[3353] = cin[2191];
assign cj_6144[3354] = cin[2358];
assign cj_6144[3355] = cin[3485];
assign cj_6144[3356] = cin[5572];
assign cj_6144[3357] = cin[2475];
assign cj_6144[3358] = cin[338];
assign cj_6144[3359] = cin[5305];
assign cj_6144[3360] = cin[5088];
assign cj_6144[3361] = cin[5831];
assign cj_6144[3362] = cin[1390];
assign cj_6144[3363] = cin[4053];
assign cj_6144[3364] = cin[1532];
assign cj_6144[3365] = cin[6115];
assign cj_6144[3366] = cin[5514];
assign cj_6144[3367] = cin[5873];
assign cj_6144[3368] = cin[1048];
assign cj_6144[3369] = cin[3327];
assign cj_6144[3370] = cin[422];
assign cj_6144[3371] = cin[4621];
assign cj_6144[3372] = cin[3636];
assign cj_6144[3373] = cin[3611];
assign cj_6144[3374] = cin[4546];
assign cj_6144[3375] = cin[297];
assign cj_6144[3376] = cin[3152];
assign cj_6144[3377] = cin[823];
assign cj_6144[3378] = cin[5598];
assign cj_6144[3379] = cin[5189];
assign cj_6144[3380] = cin[5740];
assign cj_6144[3381] = cin[1107];
assign cj_6144[3382] = cin[3578];
assign cj_6144[3383] = cin[865];
assign cj_6144[3384] = cin[5256];
assign cj_6144[3385] = cin[4463];
assign cj_6144[3386] = cin[4630];
assign cj_6144[3387] = cin[5757];
assign cj_6144[3388] = cin[1700];
assign cj_6144[3389] = cin[4747];
assign cj_6144[3390] = cin[2610];
assign cj_6144[3391] = cin[1433];
assign cj_6144[3392] = cin[1216];
assign cj_6144[3393] = cin[1959];
assign cj_6144[3394] = cin[3662];
assign cj_6144[3395] = cin[181];
assign cj_6144[3396] = cin[3804];
assign cj_6144[3397] = cin[2243];
assign cj_6144[3398] = cin[1642];
assign cj_6144[3399] = cin[2001];
assign cj_6144[3400] = cin[3320];
assign cj_6144[3401] = cin[5599];
assign cj_6144[3402] = cin[2694];
assign cj_6144[3403] = cin[749];
assign cj_6144[3404] = cin[5908];
assign cj_6144[3405] = cin[5883];
assign cj_6144[3406] = cin[674];
assign cj_6144[3407] = cin[2569];
assign cj_6144[3408] = cin[5424];
assign cj_6144[3409] = cin[3095];
assign cj_6144[3410] = cin[1726];
assign cj_6144[3411] = cin[1317];
assign cj_6144[3412] = cin[1868];
assign cj_6144[3413] = cin[3379];
assign cj_6144[3414] = cin[5850];
assign cj_6144[3415] = cin[3137];
assign cj_6144[3416] = cin[1384];
assign cj_6144[3417] = cin[591];
assign cj_6144[3418] = cin[758];
assign cj_6144[3419] = cin[1885];
assign cj_6144[3420] = cin[3972];
assign cj_6144[3421] = cin[875];
assign cj_6144[3422] = cin[4882];
assign cj_6144[3423] = cin[3705];
assign cj_6144[3424] = cin[3488];
assign cj_6144[3425] = cin[4231];
assign cj_6144[3426] = cin[5934];
assign cj_6144[3427] = cin[2453];
assign cj_6144[3428] = cin[6076];
assign cj_6144[3429] = cin[4515];
assign cj_6144[3430] = cin[3914];
assign cj_6144[3431] = cin[4273];
assign cj_6144[3432] = cin[5592];
assign cj_6144[3433] = cin[1727];
assign cj_6144[3434] = cin[4966];
assign cj_6144[3435] = cin[3021];
assign cj_6144[3436] = cin[2036];
assign cj_6144[3437] = cin[2011];
assign cj_6144[3438] = cin[2946];
assign cj_6144[3439] = cin[4841];
assign cj_6144[3440] = cin[1552];
assign cj_6144[3441] = cin[5367];
assign cj_6144[3442] = cin[3998];
assign cj_6144[3443] = cin[3589];
assign cj_6144[3444] = cin[4140];
assign cj_6144[3445] = cin[5651];
assign cj_6144[3446] = cin[1978];
assign cj_6144[3447] = cin[5409];
assign cj_6144[3448] = cin[3656];
assign cj_6144[3449] = cin[2863];
assign cj_6144[3450] = cin[3030];
assign cj_6144[3451] = cin[4157];
assign cj_6144[3452] = cin[100];
assign cj_6144[3453] = cin[3147];
assign cj_6144[3454] = cin[1010];
assign cj_6144[3455] = cin[5977];
assign cj_6144[3456] = cin[5760];
assign cj_6144[3457] = cin[359];
assign cj_6144[3458] = cin[2062];
assign cj_6144[3459] = cin[4725];
assign cj_6144[3460] = cin[2204];
assign cj_6144[3461] = cin[643];
assign cj_6144[3462] = cin[42];
assign cj_6144[3463] = cin[401];
assign cj_6144[3464] = cin[1720];
assign cj_6144[3465] = cin[3999];
assign cj_6144[3466] = cin[1094];
assign cj_6144[3467] = cin[5293];
assign cj_6144[3468] = cin[4308];
assign cj_6144[3469] = cin[4283];
assign cj_6144[3470] = cin[5218];
assign cj_6144[3471] = cin[969];
assign cj_6144[3472] = cin[3824];
assign cj_6144[3473] = cin[1495];
assign cj_6144[3474] = cin[126];
assign cj_6144[3475] = cin[5861];
assign cj_6144[3476] = cin[268];
assign cj_6144[3477] = cin[1779];
assign cj_6144[3478] = cin[4250];
assign cj_6144[3479] = cin[1537];
assign cj_6144[3480] = cin[5928];
assign cj_6144[3481] = cin[5135];
assign cj_6144[3482] = cin[5302];
assign cj_6144[3483] = cin[285];
assign cj_6144[3484] = cin[2372];
assign cj_6144[3485] = cin[5419];
assign cj_6144[3486] = cin[3282];
assign cj_6144[3487] = cin[2105];
assign cj_6144[3488] = cin[1888];
assign cj_6144[3489] = cin[2631];
assign cj_6144[3490] = cin[4334];
assign cj_6144[3491] = cin[853];
assign cj_6144[3492] = cin[4476];
assign cj_6144[3493] = cin[2915];
assign cj_6144[3494] = cin[2314];
assign cj_6144[3495] = cin[2673];
assign cj_6144[3496] = cin[3992];
assign cj_6144[3497] = cin[127];
assign cj_6144[3498] = cin[3366];
assign cj_6144[3499] = cin[1421];
assign cj_6144[3500] = cin[436];
assign cj_6144[3501] = cin[411];
assign cj_6144[3502] = cin[1346];
assign cj_6144[3503] = cin[3241];
assign cj_6144[3504] = cin[6096];
assign cj_6144[3505] = cin[3767];
assign cj_6144[3506] = cin[2398];
assign cj_6144[3507] = cin[1989];
assign cj_6144[3508] = cin[2540];
assign cj_6144[3509] = cin[4051];
assign cj_6144[3510] = cin[378];
assign cj_6144[3511] = cin[3809];
assign cj_6144[3512] = cin[2056];
assign cj_6144[3513] = cin[1263];
assign cj_6144[3514] = cin[1430];
assign cj_6144[3515] = cin[2557];
assign cj_6144[3516] = cin[4644];
assign cj_6144[3517] = cin[1547];
assign cj_6144[3518] = cin[5554];
assign cj_6144[3519] = cin[4377];
assign cj_6144[3520] = cin[4160];
assign cj_6144[3521] = cin[4903];
assign cj_6144[3522] = cin[462];
assign cj_6144[3523] = cin[3125];
assign cj_6144[3524] = cin[604];
assign cj_6144[3525] = cin[5187];
assign cj_6144[3526] = cin[4586];
assign cj_6144[3527] = cin[4945];
assign cj_6144[3528] = cin[120];
assign cj_6144[3529] = cin[2399];
assign cj_6144[3530] = cin[5638];
assign cj_6144[3531] = cin[3693];
assign cj_6144[3532] = cin[2708];
assign cj_6144[3533] = cin[2683];
assign cj_6144[3534] = cin[3618];
assign cj_6144[3535] = cin[5513];
assign cj_6144[3536] = cin[2224];
assign cj_6144[3537] = cin[6039];
assign cj_6144[3538] = cin[4670];
assign cj_6144[3539] = cin[4261];
assign cj_6144[3540] = cin[4812];
assign cj_6144[3541] = cin[179];
assign cj_6144[3542] = cin[2650];
assign cj_6144[3543] = cin[6081];
assign cj_6144[3544] = cin[4328];
assign cj_6144[3545] = cin[3535];
assign cj_6144[3546] = cin[3702];
assign cj_6144[3547] = cin[4829];
assign cj_6144[3548] = cin[772];
assign cj_6144[3549] = cin[3819];
assign cj_6144[3550] = cin[1682];
assign cj_6144[3551] = cin[505];
assign cj_6144[3552] = cin[288];
assign cj_6144[3553] = cin[1031];
assign cj_6144[3554] = cin[2734];
assign cj_6144[3555] = cin[5397];
assign cj_6144[3556] = cin[2876];
assign cj_6144[3557] = cin[1315];
assign cj_6144[3558] = cin[714];
assign cj_6144[3559] = cin[1073];
assign cj_6144[3560] = cin[2392];
assign cj_6144[3561] = cin[4671];
assign cj_6144[3562] = cin[1766];
assign cj_6144[3563] = cin[5965];
assign cj_6144[3564] = cin[4980];
assign cj_6144[3565] = cin[4955];
assign cj_6144[3566] = cin[5890];
assign cj_6144[3567] = cin[1641];
assign cj_6144[3568] = cin[4496];
assign cj_6144[3569] = cin[2167];
assign cj_6144[3570] = cin[798];
assign cj_6144[3571] = cin[389];
assign cj_6144[3572] = cin[940];
assign cj_6144[3573] = cin[2451];
assign cj_6144[3574] = cin[4922];
assign cj_6144[3575] = cin[2209];
assign cj_6144[3576] = cin[456];
assign cj_6144[3577] = cin[5807];
assign cj_6144[3578] = cin[5974];
assign cj_6144[3579] = cin[957];
assign cj_6144[3580] = cin[3044];
assign cj_6144[3581] = cin[6091];
assign cj_6144[3582] = cin[3954];
assign cj_6144[3583] = cin[2777];
assign cj_6144[3584] = cin[2560];
assign cj_6144[3585] = cin[3303];
assign cj_6144[3586] = cin[5006];
assign cj_6144[3587] = cin[1525];
assign cj_6144[3588] = cin[5148];
assign cj_6144[3589] = cin[3587];
assign cj_6144[3590] = cin[2986];
assign cj_6144[3591] = cin[3345];
assign cj_6144[3592] = cin[4664];
assign cj_6144[3593] = cin[799];
assign cj_6144[3594] = cin[4038];
assign cj_6144[3595] = cin[2093];
assign cj_6144[3596] = cin[1108];
assign cj_6144[3597] = cin[1083];
assign cj_6144[3598] = cin[2018];
assign cj_6144[3599] = cin[3913];
assign cj_6144[3600] = cin[624];
assign cj_6144[3601] = cin[4439];
assign cj_6144[3602] = cin[3070];
assign cj_6144[3603] = cin[2661];
assign cj_6144[3604] = cin[3212];
assign cj_6144[3605] = cin[4723];
assign cj_6144[3606] = cin[1050];
assign cj_6144[3607] = cin[4481];
assign cj_6144[3608] = cin[2728];
assign cj_6144[3609] = cin[1935];
assign cj_6144[3610] = cin[2102];
assign cj_6144[3611] = cin[3229];
assign cj_6144[3612] = cin[5316];
assign cj_6144[3613] = cin[2219];
assign cj_6144[3614] = cin[82];
assign cj_6144[3615] = cin[5049];
assign cj_6144[3616] = cin[4832];
assign cj_6144[3617] = cin[5575];
assign cj_6144[3618] = cin[1134];
assign cj_6144[3619] = cin[3797];
assign cj_6144[3620] = cin[1276];
assign cj_6144[3621] = cin[5859];
assign cj_6144[3622] = cin[5258];
assign cj_6144[3623] = cin[5617];
assign cj_6144[3624] = cin[792];
assign cj_6144[3625] = cin[3071];
assign cj_6144[3626] = cin[166];
assign cj_6144[3627] = cin[4365];
assign cj_6144[3628] = cin[3380];
assign cj_6144[3629] = cin[3355];
assign cj_6144[3630] = cin[4290];
assign cj_6144[3631] = cin[41];
assign cj_6144[3632] = cin[2896];
assign cj_6144[3633] = cin[567];
assign cj_6144[3634] = cin[5342];
assign cj_6144[3635] = cin[4933];
assign cj_6144[3636] = cin[5484];
assign cj_6144[3637] = cin[851];
assign cj_6144[3638] = cin[3322];
assign cj_6144[3639] = cin[609];
assign cj_6144[3640] = cin[5000];
assign cj_6144[3641] = cin[4207];
assign cj_6144[3642] = cin[4374];
assign cj_6144[3643] = cin[5501];
assign cj_6144[3644] = cin[1444];
assign cj_6144[3645] = cin[4491];
assign cj_6144[3646] = cin[2354];
assign cj_6144[3647] = cin[1177];
assign cj_6144[3648] = cin[960];
assign cj_6144[3649] = cin[1703];
assign cj_6144[3650] = cin[3406];
assign cj_6144[3651] = cin[6069];
assign cj_6144[3652] = cin[3548];
assign cj_6144[3653] = cin[1987];
assign cj_6144[3654] = cin[1386];
assign cj_6144[3655] = cin[1745];
assign cj_6144[3656] = cin[3064];
assign cj_6144[3657] = cin[5343];
assign cj_6144[3658] = cin[2438];
assign cj_6144[3659] = cin[493];
assign cj_6144[3660] = cin[5652];
assign cj_6144[3661] = cin[5627];
assign cj_6144[3662] = cin[418];
assign cj_6144[3663] = cin[2313];
assign cj_6144[3664] = cin[5168];
assign cj_6144[3665] = cin[2839];
assign cj_6144[3666] = cin[1470];
assign cj_6144[3667] = cin[1061];
assign cj_6144[3668] = cin[1612];
assign cj_6144[3669] = cin[3123];
assign cj_6144[3670] = cin[5594];
assign cj_6144[3671] = cin[2881];
assign cj_6144[3672] = cin[1128];
assign cj_6144[3673] = cin[335];
assign cj_6144[3674] = cin[502];
assign cj_6144[3675] = cin[1629];
assign cj_6144[3676] = cin[3716];
assign cj_6144[3677] = cin[619];
assign cj_6144[3678] = cin[4626];
assign cj_6144[3679] = cin[3449];
assign cj_6144[3680] = cin[3232];
assign cj_6144[3681] = cin[3975];
assign cj_6144[3682] = cin[5678];
assign cj_6144[3683] = cin[2197];
assign cj_6144[3684] = cin[5820];
assign cj_6144[3685] = cin[4259];
assign cj_6144[3686] = cin[3658];
assign cj_6144[3687] = cin[4017];
assign cj_6144[3688] = cin[5336];
assign cj_6144[3689] = cin[1471];
assign cj_6144[3690] = cin[4710];
assign cj_6144[3691] = cin[2765];
assign cj_6144[3692] = cin[1780];
assign cj_6144[3693] = cin[1755];
assign cj_6144[3694] = cin[2690];
assign cj_6144[3695] = cin[4585];
assign cj_6144[3696] = cin[1296];
assign cj_6144[3697] = cin[5111];
assign cj_6144[3698] = cin[3742];
assign cj_6144[3699] = cin[3333];
assign cj_6144[3700] = cin[3884];
assign cj_6144[3701] = cin[5395];
assign cj_6144[3702] = cin[1722];
assign cj_6144[3703] = cin[5153];
assign cj_6144[3704] = cin[3400];
assign cj_6144[3705] = cin[2607];
assign cj_6144[3706] = cin[2774];
assign cj_6144[3707] = cin[3901];
assign cj_6144[3708] = cin[5988];
assign cj_6144[3709] = cin[2891];
assign cj_6144[3710] = cin[754];
assign cj_6144[3711] = cin[5721];
assign cj_6144[3712] = cin[5504];
assign cj_6144[3713] = cin[103];
assign cj_6144[3714] = cin[1806];
assign cj_6144[3715] = cin[4469];
assign cj_6144[3716] = cin[1948];
assign cj_6144[3717] = cin[387];
assign cj_6144[3718] = cin[5930];
assign cj_6144[3719] = cin[145];
assign cj_6144[3720] = cin[1464];
assign cj_6144[3721] = cin[3743];
assign cj_6144[3722] = cin[838];
assign cj_6144[3723] = cin[5037];
assign cj_6144[3724] = cin[4052];
assign cj_6144[3725] = cin[4027];
assign cj_6144[3726] = cin[4962];
assign cj_6144[3727] = cin[713];
assign cj_6144[3728] = cin[3568];
assign cj_6144[3729] = cin[1239];
assign cj_6144[3730] = cin[6014];
assign cj_6144[3731] = cin[5605];
assign cj_6144[3732] = cin[12];
assign cj_6144[3733] = cin[1523];
assign cj_6144[3734] = cin[3994];
assign cj_6144[3735] = cin[1281];
assign cj_6144[3736] = cin[5672];
assign cj_6144[3737] = cin[4879];
assign cj_6144[3738] = cin[5046];
assign cj_6144[3739] = cin[29];
assign cj_6144[3740] = cin[2116];
assign cj_6144[3741] = cin[5163];
assign cj_6144[3742] = cin[3026];
assign cj_6144[3743] = cin[1849];
assign cj_6144[3744] = cin[1632];
assign cj_6144[3745] = cin[2375];
assign cj_6144[3746] = cin[4078];
assign cj_6144[3747] = cin[597];
assign cj_6144[3748] = cin[4220];
assign cj_6144[3749] = cin[2659];
assign cj_6144[3750] = cin[2058];
assign cj_6144[3751] = cin[2417];
assign cj_6144[3752] = cin[3736];
assign cj_6144[3753] = cin[6015];
assign cj_6144[3754] = cin[3110];
assign cj_6144[3755] = cin[1165];
assign cj_6144[3756] = cin[180];
assign cj_6144[3757] = cin[155];
assign cj_6144[3758] = cin[1090];
assign cj_6144[3759] = cin[2985];
assign cj_6144[3760] = cin[5840];
assign cj_6144[3761] = cin[3511];
assign cj_6144[3762] = cin[2142];
assign cj_6144[3763] = cin[1733];
assign cj_6144[3764] = cin[2284];
assign cj_6144[3765] = cin[3795];
assign cj_6144[3766] = cin[122];
assign cj_6144[3767] = cin[3553];
assign cj_6144[3768] = cin[1800];
assign cj_6144[3769] = cin[1007];
assign cj_6144[3770] = cin[1174];
assign cj_6144[3771] = cin[2301];
assign cj_6144[3772] = cin[4388];
assign cj_6144[3773] = cin[1291];
assign cj_6144[3774] = cin[5298];
assign cj_6144[3775] = cin[4121];
assign cj_6144[3776] = cin[3904];
assign cj_6144[3777] = cin[4647];
assign cj_6144[3778] = cin[206];
assign cj_6144[3779] = cin[2869];
assign cj_6144[3780] = cin[348];
assign cj_6144[3781] = cin[4931];
assign cj_6144[3782] = cin[4330];
assign cj_6144[3783] = cin[4689];
assign cj_6144[3784] = cin[6008];
assign cj_6144[3785] = cin[2143];
assign cj_6144[3786] = cin[5382];
assign cj_6144[3787] = cin[3437];
assign cj_6144[3788] = cin[2452];
assign cj_6144[3789] = cin[2427];
assign cj_6144[3790] = cin[3362];
assign cj_6144[3791] = cin[5257];
assign cj_6144[3792] = cin[1968];
assign cj_6144[3793] = cin[5783];
assign cj_6144[3794] = cin[4414];
assign cj_6144[3795] = cin[4005];
assign cj_6144[3796] = cin[4556];
assign cj_6144[3797] = cin[6067];
assign cj_6144[3798] = cin[2394];
assign cj_6144[3799] = cin[5825];
assign cj_6144[3800] = cin[4072];
assign cj_6144[3801] = cin[3279];
assign cj_6144[3802] = cin[3446];
assign cj_6144[3803] = cin[4573];
assign cj_6144[3804] = cin[516];
assign cj_6144[3805] = cin[3563];
assign cj_6144[3806] = cin[1426];
assign cj_6144[3807] = cin[249];
assign cj_6144[3808] = cin[32];
assign cj_6144[3809] = cin[775];
assign cj_6144[3810] = cin[2478];
assign cj_6144[3811] = cin[5141];
assign cj_6144[3812] = cin[2620];
assign cj_6144[3813] = cin[1059];
assign cj_6144[3814] = cin[458];
assign cj_6144[3815] = cin[817];
assign cj_6144[3816] = cin[2136];
assign cj_6144[3817] = cin[4415];
assign cj_6144[3818] = cin[1510];
assign cj_6144[3819] = cin[5709];
assign cj_6144[3820] = cin[4724];
assign cj_6144[3821] = cin[4699];
assign cj_6144[3822] = cin[5634];
assign cj_6144[3823] = cin[1385];
assign cj_6144[3824] = cin[4240];
assign cj_6144[3825] = cin[1911];
assign cj_6144[3826] = cin[542];
assign cj_6144[3827] = cin[133];
assign cj_6144[3828] = cin[684];
assign cj_6144[3829] = cin[2195];
assign cj_6144[3830] = cin[4666];
assign cj_6144[3831] = cin[1953];
assign cj_6144[3832] = cin[200];
assign cj_6144[3833] = cin[5551];
assign cj_6144[3834] = cin[5718];
assign cj_6144[3835] = cin[701];
assign cj_6144[3836] = cin[2788];
assign cj_6144[3837] = cin[5835];
assign cj_6144[3838] = cin[3698];
assign cj_6144[3839] = cin[2521];
assign cj_6144[3840] = cin[2304];
assign cj_6144[3841] = cin[3047];
assign cj_6144[3842] = cin[4750];
assign cj_6144[3843] = cin[1269];
assign cj_6144[3844] = cin[4892];
assign cj_6144[3845] = cin[3331];
assign cj_6144[3846] = cin[2730];
assign cj_6144[3847] = cin[3089];
assign cj_6144[3848] = cin[4408];
assign cj_6144[3849] = cin[543];
assign cj_6144[3850] = cin[3782];
assign cj_6144[3851] = cin[1837];
assign cj_6144[3852] = cin[852];
assign cj_6144[3853] = cin[827];
assign cj_6144[3854] = cin[1762];
assign cj_6144[3855] = cin[3657];
assign cj_6144[3856] = cin[368];
assign cj_6144[3857] = cin[4183];
assign cj_6144[3858] = cin[2814];
assign cj_6144[3859] = cin[2405];
assign cj_6144[3860] = cin[2956];
assign cj_6144[3861] = cin[4467];
assign cj_6144[3862] = cin[794];
assign cj_6144[3863] = cin[4225];
assign cj_6144[3864] = cin[2472];
assign cj_6144[3865] = cin[1679];
assign cj_6144[3866] = cin[1846];
assign cj_6144[3867] = cin[2973];
assign cj_6144[3868] = cin[5060];
assign cj_6144[3869] = cin[1963];
assign cj_6144[3870] = cin[5970];
assign cj_6144[3871] = cin[4793];
assign cj_6144[3872] = cin[4576];
assign cj_6144[3873] = cin[5319];
assign cj_6144[3874] = cin[878];
assign cj_6144[3875] = cin[3541];
assign cj_6144[3876] = cin[1020];
assign cj_6144[3877] = cin[5603];
assign cj_6144[3878] = cin[5002];
assign cj_6144[3879] = cin[5361];
assign cj_6144[3880] = cin[536];
assign cj_6144[3881] = cin[2815];
assign cj_6144[3882] = cin[6054];
assign cj_6144[3883] = cin[4109];
assign cj_6144[3884] = cin[3124];
assign cj_6144[3885] = cin[3099];
assign cj_6144[3886] = cin[4034];
assign cj_6144[3887] = cin[5929];
assign cj_6144[3888] = cin[2640];
assign cj_6144[3889] = cin[311];
assign cj_6144[3890] = cin[5086];
assign cj_6144[3891] = cin[4677];
assign cj_6144[3892] = cin[5228];
assign cj_6144[3893] = cin[595];
assign cj_6144[3894] = cin[3066];
assign cj_6144[3895] = cin[353];
assign cj_6144[3896] = cin[4744];
assign cj_6144[3897] = cin[3951];
assign cj_6144[3898] = cin[4118];
assign cj_6144[3899] = cin[5245];
assign cj_6144[3900] = cin[1188];
assign cj_6144[3901] = cin[4235];
assign cj_6144[3902] = cin[2098];
assign cj_6144[3903] = cin[921];
assign cj_6144[3904] = cin[704];
assign cj_6144[3905] = cin[1447];
assign cj_6144[3906] = cin[3150];
assign cj_6144[3907] = cin[5813];
assign cj_6144[3908] = cin[3292];
assign cj_6144[3909] = cin[1731];
assign cj_6144[3910] = cin[1130];
assign cj_6144[3911] = cin[1489];
assign cj_6144[3912] = cin[2808];
assign cj_6144[3913] = cin[5087];
assign cj_6144[3914] = cin[2182];
assign cj_6144[3915] = cin[237];
assign cj_6144[3916] = cin[5396];
assign cj_6144[3917] = cin[5371];
assign cj_6144[3918] = cin[162];
assign cj_6144[3919] = cin[2057];
assign cj_6144[3920] = cin[4912];
assign cj_6144[3921] = cin[2583];
assign cj_6144[3922] = cin[1214];
assign cj_6144[3923] = cin[805];
assign cj_6144[3924] = cin[1356];
assign cj_6144[3925] = cin[2867];
assign cj_6144[3926] = cin[5338];
assign cj_6144[3927] = cin[2625];
assign cj_6144[3928] = cin[872];
assign cj_6144[3929] = cin[79];
assign cj_6144[3930] = cin[246];
assign cj_6144[3931] = cin[1373];
assign cj_6144[3932] = cin[3460];
assign cj_6144[3933] = cin[363];
assign cj_6144[3934] = cin[4370];
assign cj_6144[3935] = cin[3193];
assign cj_6144[3936] = cin[2976];
assign cj_6144[3937] = cin[3719];
assign cj_6144[3938] = cin[5422];
assign cj_6144[3939] = cin[1941];
assign cj_6144[3940] = cin[5564];
assign cj_6144[3941] = cin[4003];
assign cj_6144[3942] = cin[3402];
assign cj_6144[3943] = cin[3761];
assign cj_6144[3944] = cin[5080];
assign cj_6144[3945] = cin[1215];
assign cj_6144[3946] = cin[4454];
assign cj_6144[3947] = cin[2509];
assign cj_6144[3948] = cin[1524];
assign cj_6144[3949] = cin[1499];
assign cj_6144[3950] = cin[2434];
assign cj_6144[3951] = cin[4329];
assign cj_6144[3952] = cin[1040];
assign cj_6144[3953] = cin[4855];
assign cj_6144[3954] = cin[3486];
assign cj_6144[3955] = cin[3077];
assign cj_6144[3956] = cin[3628];
assign cj_6144[3957] = cin[5139];
assign cj_6144[3958] = cin[1466];
assign cj_6144[3959] = cin[4897];
assign cj_6144[3960] = cin[3144];
assign cj_6144[3961] = cin[2351];
assign cj_6144[3962] = cin[2518];
assign cj_6144[3963] = cin[3645];
assign cj_6144[3964] = cin[5732];
assign cj_6144[3965] = cin[2635];
assign cj_6144[3966] = cin[498];
assign cj_6144[3967] = cin[5465];
assign cj_6144[3968] = cin[5248];
assign cj_6144[3969] = cin[5991];
assign cj_6144[3970] = cin[1550];
assign cj_6144[3971] = cin[4213];
assign cj_6144[3972] = cin[1692];
assign cj_6144[3973] = cin[131];
assign cj_6144[3974] = cin[5674];
assign cj_6144[3975] = cin[6033];
assign cj_6144[3976] = cin[1208];
assign cj_6144[3977] = cin[3487];
assign cj_6144[3978] = cin[582];
assign cj_6144[3979] = cin[4781];
assign cj_6144[3980] = cin[3796];
assign cj_6144[3981] = cin[3771];
assign cj_6144[3982] = cin[4706];
assign cj_6144[3983] = cin[457];
assign cj_6144[3984] = cin[3312];
assign cj_6144[3985] = cin[983];
assign cj_6144[3986] = cin[5758];
assign cj_6144[3987] = cin[5349];
assign cj_6144[3988] = cin[5900];
assign cj_6144[3989] = cin[1267];
assign cj_6144[3990] = cin[3738];
assign cj_6144[3991] = cin[1025];
assign cj_6144[3992] = cin[5416];
assign cj_6144[3993] = cin[4623];
assign cj_6144[3994] = cin[4790];
assign cj_6144[3995] = cin[5917];
assign cj_6144[3996] = cin[1860];
assign cj_6144[3997] = cin[4907];
assign cj_6144[3998] = cin[2770];
assign cj_6144[3999] = cin[1593];
assign cj_6144[4000] = cin[1376];
assign cj_6144[4001] = cin[2119];
assign cj_6144[4002] = cin[3822];
assign cj_6144[4003] = cin[341];
assign cj_6144[4004] = cin[3964];
assign cj_6144[4005] = cin[2403];
assign cj_6144[4006] = cin[1802];
assign cj_6144[4007] = cin[2161];
assign cj_6144[4008] = cin[3480];
assign cj_6144[4009] = cin[5759];
assign cj_6144[4010] = cin[2854];
assign cj_6144[4011] = cin[909];
assign cj_6144[4012] = cin[6068];
assign cj_6144[4013] = cin[6043];
assign cj_6144[4014] = cin[834];
assign cj_6144[4015] = cin[2729];
assign cj_6144[4016] = cin[5584];
assign cj_6144[4017] = cin[3255];
assign cj_6144[4018] = cin[1886];
assign cj_6144[4019] = cin[1477];
assign cj_6144[4020] = cin[2028];
assign cj_6144[4021] = cin[3539];
assign cj_6144[4022] = cin[6010];
assign cj_6144[4023] = cin[3297];
assign cj_6144[4024] = cin[1544];
assign cj_6144[4025] = cin[751];
assign cj_6144[4026] = cin[918];
assign cj_6144[4027] = cin[2045];
assign cj_6144[4028] = cin[4132];
assign cj_6144[4029] = cin[1035];
assign cj_6144[4030] = cin[5042];
assign cj_6144[4031] = cin[3865];
assign cj_6144[4032] = cin[3648];
assign cj_6144[4033] = cin[4391];
assign cj_6144[4034] = cin[6094];
assign cj_6144[4035] = cin[2613];
assign cj_6144[4036] = cin[92];
assign cj_6144[4037] = cin[4675];
assign cj_6144[4038] = cin[4074];
assign cj_6144[4039] = cin[4433];
assign cj_6144[4040] = cin[5752];
assign cj_6144[4041] = cin[1887];
assign cj_6144[4042] = cin[5126];
assign cj_6144[4043] = cin[3181];
assign cj_6144[4044] = cin[2196];
assign cj_6144[4045] = cin[2171];
assign cj_6144[4046] = cin[3106];
assign cj_6144[4047] = cin[5001];
assign cj_6144[4048] = cin[1712];
assign cj_6144[4049] = cin[5527];
assign cj_6144[4050] = cin[4158];
assign cj_6144[4051] = cin[3749];
assign cj_6144[4052] = cin[4300];
assign cj_6144[4053] = cin[5811];
assign cj_6144[4054] = cin[2138];
assign cj_6144[4055] = cin[5569];
assign cj_6144[4056] = cin[3816];
assign cj_6144[4057] = cin[3023];
assign cj_6144[4058] = cin[3190];
assign cj_6144[4059] = cin[4317];
assign cj_6144[4060] = cin[260];
assign cj_6144[4061] = cin[3307];
assign cj_6144[4062] = cin[1170];
assign cj_6144[4063] = cin[6137];
assign cj_6144[4064] = cin[5920];
assign cj_6144[4065] = cin[519];
assign cj_6144[4066] = cin[2222];
assign cj_6144[4067] = cin[4885];
assign cj_6144[4068] = cin[2364];
assign cj_6144[4069] = cin[803];
assign cj_6144[4070] = cin[202];
assign cj_6144[4071] = cin[561];
assign cj_6144[4072] = cin[1880];
assign cj_6144[4073] = cin[4159];
assign cj_6144[4074] = cin[1254];
assign cj_6144[4075] = cin[5453];
assign cj_6144[4076] = cin[4468];
assign cj_6144[4077] = cin[4443];
assign cj_6144[4078] = cin[5378];
assign cj_6144[4079] = cin[1129];
assign cj_6144[4080] = cin[3984];
assign cj_6144[4081] = cin[1655];
assign cj_6144[4082] = cin[286];
assign cj_6144[4083] = cin[6021];
assign cj_6144[4084] = cin[428];
assign cj_6144[4085] = cin[1939];
assign cj_6144[4086] = cin[4410];
assign cj_6144[4087] = cin[1697];
assign cj_6144[4088] = cin[6088];
assign cj_6144[4089] = cin[5295];
assign cj_6144[4090] = cin[5462];
assign cj_6144[4091] = cin[445];
assign cj_6144[4092] = cin[2532];
assign cj_6144[4093] = cin[5579];
assign cj_6144[4094] = cin[3442];
assign cj_6144[4095] = cin[2265];
assign cj_6144[4096] = cin[2048];
assign cj_6144[4097] = cin[2791];
assign cj_6144[4098] = cin[4494];
assign cj_6144[4099] = cin[1013];
assign cj_6144[4100] = cin[4636];
assign cj_6144[4101] = cin[3075];
assign cj_6144[4102] = cin[2474];
assign cj_6144[4103] = cin[2833];
assign cj_6144[4104] = cin[4152];
assign cj_6144[4105] = cin[287];
assign cj_6144[4106] = cin[3526];
assign cj_6144[4107] = cin[1581];
assign cj_6144[4108] = cin[596];
assign cj_6144[4109] = cin[571];
assign cj_6144[4110] = cin[1506];
assign cj_6144[4111] = cin[3401];
assign cj_6144[4112] = cin[112];
assign cj_6144[4113] = cin[3927];
assign cj_6144[4114] = cin[2558];
assign cj_6144[4115] = cin[2149];
assign cj_6144[4116] = cin[2700];
assign cj_6144[4117] = cin[4211];
assign cj_6144[4118] = cin[538];
assign cj_6144[4119] = cin[3969];
assign cj_6144[4120] = cin[2216];
assign cj_6144[4121] = cin[1423];
assign cj_6144[4122] = cin[1590];
assign cj_6144[4123] = cin[2717];
assign cj_6144[4124] = cin[4804];
assign cj_6144[4125] = cin[1707];
assign cj_6144[4126] = cin[5714];
assign cj_6144[4127] = cin[4537];
assign cj_6144[4128] = cin[4320];
assign cj_6144[4129] = cin[5063];
assign cj_6144[4130] = cin[622];
assign cj_6144[4131] = cin[3285];
assign cj_6144[4132] = cin[764];
assign cj_6144[4133] = cin[5347];
assign cj_6144[4134] = cin[4746];
assign cj_6144[4135] = cin[5105];
assign cj_6144[4136] = cin[280];
assign cj_6144[4137] = cin[2559];
assign cj_6144[4138] = cin[5798];
assign cj_6144[4139] = cin[3853];
assign cj_6144[4140] = cin[2868];
assign cj_6144[4141] = cin[2843];
assign cj_6144[4142] = cin[3778];
assign cj_6144[4143] = cin[5673];
assign cj_6144[4144] = cin[2384];
assign cj_6144[4145] = cin[55];
assign cj_6144[4146] = cin[4830];
assign cj_6144[4147] = cin[4421];
assign cj_6144[4148] = cin[4972];
assign cj_6144[4149] = cin[339];
assign cj_6144[4150] = cin[2810];
assign cj_6144[4151] = cin[97];
assign cj_6144[4152] = cin[4488];
assign cj_6144[4153] = cin[3695];
assign cj_6144[4154] = cin[3862];
assign cj_6144[4155] = cin[4989];
assign cj_6144[4156] = cin[932];
assign cj_6144[4157] = cin[3979];
assign cj_6144[4158] = cin[1842];
assign cj_6144[4159] = cin[665];
assign cj_6144[4160] = cin[448];
assign cj_6144[4161] = cin[1191];
assign cj_6144[4162] = cin[2894];
assign cj_6144[4163] = cin[5557];
assign cj_6144[4164] = cin[3036];
assign cj_6144[4165] = cin[1475];
assign cj_6144[4166] = cin[874];
assign cj_6144[4167] = cin[1233];
assign cj_6144[4168] = cin[2552];
assign cj_6144[4169] = cin[4831];
assign cj_6144[4170] = cin[1926];
assign cj_6144[4171] = cin[6125];
assign cj_6144[4172] = cin[5140];
assign cj_6144[4173] = cin[5115];
assign cj_6144[4174] = cin[6050];
assign cj_6144[4175] = cin[1801];
assign cj_6144[4176] = cin[4656];
assign cj_6144[4177] = cin[2327];
assign cj_6144[4178] = cin[958];
assign cj_6144[4179] = cin[549];
assign cj_6144[4180] = cin[1100];
assign cj_6144[4181] = cin[2611];
assign cj_6144[4182] = cin[5082];
assign cj_6144[4183] = cin[2369];
assign cj_6144[4184] = cin[616];
assign cj_6144[4185] = cin[5967];
assign cj_6144[4186] = cin[6134];
assign cj_6144[4187] = cin[1117];
assign cj_6144[4188] = cin[3204];
assign cj_6144[4189] = cin[107];
assign cj_6144[4190] = cin[4114];
assign cj_6144[4191] = cin[2937];
assign cj_6144[4192] = cin[2720];
assign cj_6144[4193] = cin[3463];
assign cj_6144[4194] = cin[5166];
assign cj_6144[4195] = cin[1685];
assign cj_6144[4196] = cin[5308];
assign cj_6144[4197] = cin[3747];
assign cj_6144[4198] = cin[3146];
assign cj_6144[4199] = cin[3505];
assign cj_6144[4200] = cin[4824];
assign cj_6144[4201] = cin[959];
assign cj_6144[4202] = cin[4198];
assign cj_6144[4203] = cin[2253];
assign cj_6144[4204] = cin[1268];
assign cj_6144[4205] = cin[1243];
assign cj_6144[4206] = cin[2178];
assign cj_6144[4207] = cin[4073];
assign cj_6144[4208] = cin[784];
assign cj_6144[4209] = cin[4599];
assign cj_6144[4210] = cin[3230];
assign cj_6144[4211] = cin[2821];
assign cj_6144[4212] = cin[3372];
assign cj_6144[4213] = cin[4883];
assign cj_6144[4214] = cin[1210];
assign cj_6144[4215] = cin[4641];
assign cj_6144[4216] = cin[2888];
assign cj_6144[4217] = cin[2095];
assign cj_6144[4218] = cin[2262];
assign cj_6144[4219] = cin[3389];
assign cj_6144[4220] = cin[5476];
assign cj_6144[4221] = cin[2379];
assign cj_6144[4222] = cin[242];
assign cj_6144[4223] = cin[5209];
assign cj_6144[4224] = cin[4992];
assign cj_6144[4225] = cin[5735];
assign cj_6144[4226] = cin[1294];
assign cj_6144[4227] = cin[3957];
assign cj_6144[4228] = cin[1436];
assign cj_6144[4229] = cin[6019];
assign cj_6144[4230] = cin[5418];
assign cj_6144[4231] = cin[5777];
assign cj_6144[4232] = cin[952];
assign cj_6144[4233] = cin[3231];
assign cj_6144[4234] = cin[326];
assign cj_6144[4235] = cin[4525];
assign cj_6144[4236] = cin[3540];
assign cj_6144[4237] = cin[3515];
assign cj_6144[4238] = cin[4450];
assign cj_6144[4239] = cin[201];
assign cj_6144[4240] = cin[3056];
assign cj_6144[4241] = cin[727];
assign cj_6144[4242] = cin[5502];
assign cj_6144[4243] = cin[5093];
assign cj_6144[4244] = cin[5644];
assign cj_6144[4245] = cin[1011];
assign cj_6144[4246] = cin[3482];
assign cj_6144[4247] = cin[769];
assign cj_6144[4248] = cin[5160];
assign cj_6144[4249] = cin[4367];
assign cj_6144[4250] = cin[4534];
assign cj_6144[4251] = cin[5661];
assign cj_6144[4252] = cin[1604];
assign cj_6144[4253] = cin[4651];
assign cj_6144[4254] = cin[2514];
assign cj_6144[4255] = cin[1337];
assign cj_6144[4256] = cin[1120];
assign cj_6144[4257] = cin[1863];
assign cj_6144[4258] = cin[3566];
assign cj_6144[4259] = cin[85];
assign cj_6144[4260] = cin[3708];
assign cj_6144[4261] = cin[2147];
assign cj_6144[4262] = cin[1546];
assign cj_6144[4263] = cin[1905];
assign cj_6144[4264] = cin[3224];
assign cj_6144[4265] = cin[5503];
assign cj_6144[4266] = cin[2598];
assign cj_6144[4267] = cin[653];
assign cj_6144[4268] = cin[5812];
assign cj_6144[4269] = cin[5787];
assign cj_6144[4270] = cin[578];
assign cj_6144[4271] = cin[2473];
assign cj_6144[4272] = cin[5328];
assign cj_6144[4273] = cin[2999];
assign cj_6144[4274] = cin[1630];
assign cj_6144[4275] = cin[1221];
assign cj_6144[4276] = cin[1772];
assign cj_6144[4277] = cin[3283];
assign cj_6144[4278] = cin[5754];
assign cj_6144[4279] = cin[3041];
assign cj_6144[4280] = cin[1288];
assign cj_6144[4281] = cin[495];
assign cj_6144[4282] = cin[662];
assign cj_6144[4283] = cin[1789];
assign cj_6144[4284] = cin[3876];
assign cj_6144[4285] = cin[779];
assign cj_6144[4286] = cin[4786];
assign cj_6144[4287] = cin[3609];
assign cj_6144[4288] = cin[3392];
assign cj_6144[4289] = cin[4135];
assign cj_6144[4290] = cin[5838];
assign cj_6144[4291] = cin[2357];
assign cj_6144[4292] = cin[5980];
assign cj_6144[4293] = cin[4419];
assign cj_6144[4294] = cin[3818];
assign cj_6144[4295] = cin[4177];
assign cj_6144[4296] = cin[5496];
assign cj_6144[4297] = cin[1631];
assign cj_6144[4298] = cin[4870];
assign cj_6144[4299] = cin[2925];
assign cj_6144[4300] = cin[1940];
assign cj_6144[4301] = cin[1915];
assign cj_6144[4302] = cin[2850];
assign cj_6144[4303] = cin[4745];
assign cj_6144[4304] = cin[1456];
assign cj_6144[4305] = cin[5271];
assign cj_6144[4306] = cin[3902];
assign cj_6144[4307] = cin[3493];
assign cj_6144[4308] = cin[4044];
assign cj_6144[4309] = cin[5555];
assign cj_6144[4310] = cin[1882];
assign cj_6144[4311] = cin[5313];
assign cj_6144[4312] = cin[3560];
assign cj_6144[4313] = cin[2767];
assign cj_6144[4314] = cin[2934];
assign cj_6144[4315] = cin[4061];
assign cj_6144[4316] = cin[4];
assign cj_6144[4317] = cin[3051];
assign cj_6144[4318] = cin[914];
assign cj_6144[4319] = cin[5881];
assign cj_6144[4320] = cin[5664];
assign cj_6144[4321] = cin[263];
assign cj_6144[4322] = cin[1966];
assign cj_6144[4323] = cin[4629];
assign cj_6144[4324] = cin[2108];
assign cj_6144[4325] = cin[547];
assign cj_6144[4326] = cin[6090];
assign cj_6144[4327] = cin[305];
assign cj_6144[4328] = cin[1624];
assign cj_6144[4329] = cin[3903];
assign cj_6144[4330] = cin[998];
assign cj_6144[4331] = cin[5197];
assign cj_6144[4332] = cin[4212];
assign cj_6144[4333] = cin[4187];
assign cj_6144[4334] = cin[5122];
assign cj_6144[4335] = cin[873];
assign cj_6144[4336] = cin[3728];
assign cj_6144[4337] = cin[1399];
assign cj_6144[4338] = cin[30];
assign cj_6144[4339] = cin[5765];
assign cj_6144[4340] = cin[172];
assign cj_6144[4341] = cin[1683];
assign cj_6144[4342] = cin[4154];
assign cj_6144[4343] = cin[1441];
assign cj_6144[4344] = cin[5832];
assign cj_6144[4345] = cin[5039];
assign cj_6144[4346] = cin[5206];
assign cj_6144[4347] = cin[189];
assign cj_6144[4348] = cin[2276];
assign cj_6144[4349] = cin[5323];
assign cj_6144[4350] = cin[3186];
assign cj_6144[4351] = cin[2009];
assign cj_6144[4352] = cin[1792];
assign cj_6144[4353] = cin[2535];
assign cj_6144[4354] = cin[4238];
assign cj_6144[4355] = cin[757];
assign cj_6144[4356] = cin[4380];
assign cj_6144[4357] = cin[2819];
assign cj_6144[4358] = cin[2218];
assign cj_6144[4359] = cin[2577];
assign cj_6144[4360] = cin[3896];
assign cj_6144[4361] = cin[31];
assign cj_6144[4362] = cin[3270];
assign cj_6144[4363] = cin[1325];
assign cj_6144[4364] = cin[340];
assign cj_6144[4365] = cin[315];
assign cj_6144[4366] = cin[1250];
assign cj_6144[4367] = cin[3145];
assign cj_6144[4368] = cin[6000];
assign cj_6144[4369] = cin[3671];
assign cj_6144[4370] = cin[2302];
assign cj_6144[4371] = cin[1893];
assign cj_6144[4372] = cin[2444];
assign cj_6144[4373] = cin[3955];
assign cj_6144[4374] = cin[282];
assign cj_6144[4375] = cin[3713];
assign cj_6144[4376] = cin[1960];
assign cj_6144[4377] = cin[1167];
assign cj_6144[4378] = cin[1334];
assign cj_6144[4379] = cin[2461];
assign cj_6144[4380] = cin[4548];
assign cj_6144[4381] = cin[1451];
assign cj_6144[4382] = cin[5458];
assign cj_6144[4383] = cin[4281];
assign cj_6144[4384] = cin[4064];
assign cj_6144[4385] = cin[4807];
assign cj_6144[4386] = cin[366];
assign cj_6144[4387] = cin[3029];
assign cj_6144[4388] = cin[508];
assign cj_6144[4389] = cin[5091];
assign cj_6144[4390] = cin[4490];
assign cj_6144[4391] = cin[4849];
assign cj_6144[4392] = cin[24];
assign cj_6144[4393] = cin[2303];
assign cj_6144[4394] = cin[5542];
assign cj_6144[4395] = cin[3597];
assign cj_6144[4396] = cin[2612];
assign cj_6144[4397] = cin[2587];
assign cj_6144[4398] = cin[3522];
assign cj_6144[4399] = cin[5417];
assign cj_6144[4400] = cin[2128];
assign cj_6144[4401] = cin[5943];
assign cj_6144[4402] = cin[4574];
assign cj_6144[4403] = cin[4165];
assign cj_6144[4404] = cin[4716];
assign cj_6144[4405] = cin[83];
assign cj_6144[4406] = cin[2554];
assign cj_6144[4407] = cin[5985];
assign cj_6144[4408] = cin[4232];
assign cj_6144[4409] = cin[3439];
assign cj_6144[4410] = cin[3606];
assign cj_6144[4411] = cin[4733];
assign cj_6144[4412] = cin[676];
assign cj_6144[4413] = cin[3723];
assign cj_6144[4414] = cin[1586];
assign cj_6144[4415] = cin[409];
assign cj_6144[4416] = cin[192];
assign cj_6144[4417] = cin[935];
assign cj_6144[4418] = cin[2638];
assign cj_6144[4419] = cin[5301];
assign cj_6144[4420] = cin[2780];
assign cj_6144[4421] = cin[1219];
assign cj_6144[4422] = cin[618];
assign cj_6144[4423] = cin[977];
assign cj_6144[4424] = cin[2296];
assign cj_6144[4425] = cin[4575];
assign cj_6144[4426] = cin[1670];
assign cj_6144[4427] = cin[5869];
assign cj_6144[4428] = cin[4884];
assign cj_6144[4429] = cin[4859];
assign cj_6144[4430] = cin[5794];
assign cj_6144[4431] = cin[1545];
assign cj_6144[4432] = cin[4400];
assign cj_6144[4433] = cin[2071];
assign cj_6144[4434] = cin[702];
assign cj_6144[4435] = cin[293];
assign cj_6144[4436] = cin[844];
assign cj_6144[4437] = cin[2355];
assign cj_6144[4438] = cin[4826];
assign cj_6144[4439] = cin[2113];
assign cj_6144[4440] = cin[360];
assign cj_6144[4441] = cin[5711];
assign cj_6144[4442] = cin[5878];
assign cj_6144[4443] = cin[861];
assign cj_6144[4444] = cin[2948];
assign cj_6144[4445] = cin[5995];
assign cj_6144[4446] = cin[3858];
assign cj_6144[4447] = cin[2681];
assign cj_6144[4448] = cin[2464];
assign cj_6144[4449] = cin[3207];
assign cj_6144[4450] = cin[4910];
assign cj_6144[4451] = cin[1429];
assign cj_6144[4452] = cin[5052];
assign cj_6144[4453] = cin[3491];
assign cj_6144[4454] = cin[2890];
assign cj_6144[4455] = cin[3249];
assign cj_6144[4456] = cin[4568];
assign cj_6144[4457] = cin[703];
assign cj_6144[4458] = cin[3942];
assign cj_6144[4459] = cin[1997];
assign cj_6144[4460] = cin[1012];
assign cj_6144[4461] = cin[987];
assign cj_6144[4462] = cin[1922];
assign cj_6144[4463] = cin[3817];
assign cj_6144[4464] = cin[528];
assign cj_6144[4465] = cin[4343];
assign cj_6144[4466] = cin[2974];
assign cj_6144[4467] = cin[2565];
assign cj_6144[4468] = cin[3116];
assign cj_6144[4469] = cin[4627];
assign cj_6144[4470] = cin[954];
assign cj_6144[4471] = cin[4385];
assign cj_6144[4472] = cin[2632];
assign cj_6144[4473] = cin[1839];
assign cj_6144[4474] = cin[2006];
assign cj_6144[4475] = cin[3133];
assign cj_6144[4476] = cin[5220];
assign cj_6144[4477] = cin[2123];
assign cj_6144[4478] = cin[6130];
assign cj_6144[4479] = cin[4953];
assign cj_6144[4480] = cin[4736];
assign cj_6144[4481] = cin[5479];
assign cj_6144[4482] = cin[1038];
assign cj_6144[4483] = cin[3701];
assign cj_6144[4484] = cin[1180];
assign cj_6144[4485] = cin[5763];
assign cj_6144[4486] = cin[5162];
assign cj_6144[4487] = cin[5521];
assign cj_6144[4488] = cin[696];
assign cj_6144[4489] = cin[2975];
assign cj_6144[4490] = cin[70];
assign cj_6144[4491] = cin[4269];
assign cj_6144[4492] = cin[3284];
assign cj_6144[4493] = cin[3259];
assign cj_6144[4494] = cin[4194];
assign cj_6144[4495] = cin[6089];
assign cj_6144[4496] = cin[2800];
assign cj_6144[4497] = cin[471];
assign cj_6144[4498] = cin[5246];
assign cj_6144[4499] = cin[4837];
assign cj_6144[4500] = cin[5388];
assign cj_6144[4501] = cin[755];
assign cj_6144[4502] = cin[3226];
assign cj_6144[4503] = cin[513];
assign cj_6144[4504] = cin[4904];
assign cj_6144[4505] = cin[4111];
assign cj_6144[4506] = cin[4278];
assign cj_6144[4507] = cin[5405];
assign cj_6144[4508] = cin[1348];
assign cj_6144[4509] = cin[4395];
assign cj_6144[4510] = cin[2258];
assign cj_6144[4511] = cin[1081];
assign cj_6144[4512] = cin[864];
assign cj_6144[4513] = cin[1607];
assign cj_6144[4514] = cin[3310];
assign cj_6144[4515] = cin[5973];
assign cj_6144[4516] = cin[3452];
assign cj_6144[4517] = cin[1891];
assign cj_6144[4518] = cin[1290];
assign cj_6144[4519] = cin[1649];
assign cj_6144[4520] = cin[2968];
assign cj_6144[4521] = cin[5247];
assign cj_6144[4522] = cin[2342];
assign cj_6144[4523] = cin[397];
assign cj_6144[4524] = cin[5556];
assign cj_6144[4525] = cin[5531];
assign cj_6144[4526] = cin[322];
assign cj_6144[4527] = cin[2217];
assign cj_6144[4528] = cin[5072];
assign cj_6144[4529] = cin[2743];
assign cj_6144[4530] = cin[1374];
assign cj_6144[4531] = cin[965];
assign cj_6144[4532] = cin[1516];
assign cj_6144[4533] = cin[3027];
assign cj_6144[4534] = cin[5498];
assign cj_6144[4535] = cin[2785];
assign cj_6144[4536] = cin[1032];
assign cj_6144[4537] = cin[239];
assign cj_6144[4538] = cin[406];
assign cj_6144[4539] = cin[1533];
assign cj_6144[4540] = cin[3620];
assign cj_6144[4541] = cin[523];
assign cj_6144[4542] = cin[4530];
assign cj_6144[4543] = cin[3353];
assign cj_6144[4544] = cin[3136];
assign cj_6144[4545] = cin[3879];
assign cj_6144[4546] = cin[5582];
assign cj_6144[4547] = cin[2101];
assign cj_6144[4548] = cin[5724];
assign cj_6144[4549] = cin[4163];
assign cj_6144[4550] = cin[3562];
assign cj_6144[4551] = cin[3921];
assign cj_6144[4552] = cin[5240];
assign cj_6144[4553] = cin[1375];
assign cj_6144[4554] = cin[4614];
assign cj_6144[4555] = cin[2669];
assign cj_6144[4556] = cin[1684];
assign cj_6144[4557] = cin[1659];
assign cj_6144[4558] = cin[2594];
assign cj_6144[4559] = cin[4489];
assign cj_6144[4560] = cin[1200];
assign cj_6144[4561] = cin[5015];
assign cj_6144[4562] = cin[3646];
assign cj_6144[4563] = cin[3237];
assign cj_6144[4564] = cin[3788];
assign cj_6144[4565] = cin[5299];
assign cj_6144[4566] = cin[1626];
assign cj_6144[4567] = cin[5057];
assign cj_6144[4568] = cin[3304];
assign cj_6144[4569] = cin[2511];
assign cj_6144[4570] = cin[2678];
assign cj_6144[4571] = cin[3805];
assign cj_6144[4572] = cin[5892];
assign cj_6144[4573] = cin[2795];
assign cj_6144[4574] = cin[658];
assign cj_6144[4575] = cin[5625];
assign cj_6144[4576] = cin[5408];
assign cj_6144[4577] = cin[7];
assign cj_6144[4578] = cin[1710];
assign cj_6144[4579] = cin[4373];
assign cj_6144[4580] = cin[1852];
assign cj_6144[4581] = cin[291];
assign cj_6144[4582] = cin[5834];
assign cj_6144[4583] = cin[49];
assign cj_6144[4584] = cin[1368];
assign cj_6144[4585] = cin[3647];
assign cj_6144[4586] = cin[742];
assign cj_6144[4587] = cin[4941];
assign cj_6144[4588] = cin[3956];
assign cj_6144[4589] = cin[3931];
assign cj_6144[4590] = cin[4866];
assign cj_6144[4591] = cin[617];
assign cj_6144[4592] = cin[3472];
assign cj_6144[4593] = cin[1143];
assign cj_6144[4594] = cin[5918];
assign cj_6144[4595] = cin[5509];
assign cj_6144[4596] = cin[6060];
assign cj_6144[4597] = cin[1427];
assign cj_6144[4598] = cin[3898];
assign cj_6144[4599] = cin[1185];
assign cj_6144[4600] = cin[5576];
assign cj_6144[4601] = cin[4783];
assign cj_6144[4602] = cin[4950];
assign cj_6144[4603] = cin[6077];
assign cj_6144[4604] = cin[2020];
assign cj_6144[4605] = cin[5067];
assign cj_6144[4606] = cin[2930];
assign cj_6144[4607] = cin[1753];
assign cj_6144[4608] = cin[1536];
assign cj_6144[4609] = cin[2279];
assign cj_6144[4610] = cin[3982];
assign cj_6144[4611] = cin[501];
assign cj_6144[4612] = cin[4124];
assign cj_6144[4613] = cin[2563];
assign cj_6144[4614] = cin[1962];
assign cj_6144[4615] = cin[2321];
assign cj_6144[4616] = cin[3640];
assign cj_6144[4617] = cin[5919];
assign cj_6144[4618] = cin[3014];
assign cj_6144[4619] = cin[1069];
assign cj_6144[4620] = cin[84];
assign cj_6144[4621] = cin[59];
assign cj_6144[4622] = cin[994];
assign cj_6144[4623] = cin[2889];
assign cj_6144[4624] = cin[5744];
assign cj_6144[4625] = cin[3415];
assign cj_6144[4626] = cin[2046];
assign cj_6144[4627] = cin[1637];
assign cj_6144[4628] = cin[2188];
assign cj_6144[4629] = cin[3699];
assign cj_6144[4630] = cin[26];
assign cj_6144[4631] = cin[3457];
assign cj_6144[4632] = cin[1704];
assign cj_6144[4633] = cin[911];
assign cj_6144[4634] = cin[1078];
assign cj_6144[4635] = cin[2205];
assign cj_6144[4636] = cin[4292];
assign cj_6144[4637] = cin[1195];
assign cj_6144[4638] = cin[5202];
assign cj_6144[4639] = cin[4025];
assign cj_6144[4640] = cin[3808];
assign cj_6144[4641] = cin[4551];
assign cj_6144[4642] = cin[110];
assign cj_6144[4643] = cin[2773];
assign cj_6144[4644] = cin[252];
assign cj_6144[4645] = cin[4835];
assign cj_6144[4646] = cin[4234];
assign cj_6144[4647] = cin[4593];
assign cj_6144[4648] = cin[5912];
assign cj_6144[4649] = cin[2047];
assign cj_6144[4650] = cin[5286];
assign cj_6144[4651] = cin[3341];
assign cj_6144[4652] = cin[2356];
assign cj_6144[4653] = cin[2331];
assign cj_6144[4654] = cin[3266];
assign cj_6144[4655] = cin[5161];
assign cj_6144[4656] = cin[1872];
assign cj_6144[4657] = cin[5687];
assign cj_6144[4658] = cin[4318];
assign cj_6144[4659] = cin[3909];
assign cj_6144[4660] = cin[4460];
assign cj_6144[4661] = cin[5971];
assign cj_6144[4662] = cin[2298];
assign cj_6144[4663] = cin[5729];
assign cj_6144[4664] = cin[3976];
assign cj_6144[4665] = cin[3183];
assign cj_6144[4666] = cin[3350];
assign cj_6144[4667] = cin[4477];
assign cj_6144[4668] = cin[420];
assign cj_6144[4669] = cin[3467];
assign cj_6144[4670] = cin[1330];
assign cj_6144[4671] = cin[153];
assign cj_6144[4672] = cin[6080];
assign cj_6144[4673] = cin[679];
assign cj_6144[4674] = cin[2382];
assign cj_6144[4675] = cin[5045];
assign cj_6144[4676] = cin[2524];
assign cj_6144[4677] = cin[963];
assign cj_6144[4678] = cin[362];
assign cj_6144[4679] = cin[721];
assign cj_6144[4680] = cin[2040];
assign cj_6144[4681] = cin[4319];
assign cj_6144[4682] = cin[1414];
assign cj_6144[4683] = cin[5613];
assign cj_6144[4684] = cin[4628];
assign cj_6144[4685] = cin[4603];
assign cj_6144[4686] = cin[5538];
assign cj_6144[4687] = cin[1289];
assign cj_6144[4688] = cin[4144];
assign cj_6144[4689] = cin[1815];
assign cj_6144[4690] = cin[446];
assign cj_6144[4691] = cin[37];
assign cj_6144[4692] = cin[588];
assign cj_6144[4693] = cin[2099];
assign cj_6144[4694] = cin[4570];
assign cj_6144[4695] = cin[1857];
assign cj_6144[4696] = cin[104];
assign cj_6144[4697] = cin[5455];
assign cj_6144[4698] = cin[5622];
assign cj_6144[4699] = cin[605];
assign cj_6144[4700] = cin[2692];
assign cj_6144[4701] = cin[5739];
assign cj_6144[4702] = cin[3602];
assign cj_6144[4703] = cin[2425];
assign cj_6144[4704] = cin[2208];
assign cj_6144[4705] = cin[2951];
assign cj_6144[4706] = cin[4654];
assign cj_6144[4707] = cin[1173];
assign cj_6144[4708] = cin[4796];
assign cj_6144[4709] = cin[3235];
assign cj_6144[4710] = cin[2634];
assign cj_6144[4711] = cin[2993];
assign cj_6144[4712] = cin[4312];
assign cj_6144[4713] = cin[447];
assign cj_6144[4714] = cin[3686];
assign cj_6144[4715] = cin[1741];
assign cj_6144[4716] = cin[756];
assign cj_6144[4717] = cin[731];
assign cj_6144[4718] = cin[1666];
assign cj_6144[4719] = cin[3561];
assign cj_6144[4720] = cin[272];
assign cj_6144[4721] = cin[4087];
assign cj_6144[4722] = cin[2718];
assign cj_6144[4723] = cin[2309];
assign cj_6144[4724] = cin[2860];
assign cj_6144[4725] = cin[4371];
assign cj_6144[4726] = cin[698];
assign cj_6144[4727] = cin[4129];
assign cj_6144[4728] = cin[2376];
assign cj_6144[4729] = cin[1583];
assign cj_6144[4730] = cin[1750];
assign cj_6144[4731] = cin[2877];
assign cj_6144[4732] = cin[4964];
assign cj_6144[4733] = cin[1867];
assign cj_6144[4734] = cin[5874];
assign cj_6144[4735] = cin[4697];
assign cj_6144[4736] = cin[4480];
assign cj_6144[4737] = cin[5223];
assign cj_6144[4738] = cin[782];
assign cj_6144[4739] = cin[3445];
assign cj_6144[4740] = cin[924];
assign cj_6144[4741] = cin[5507];
assign cj_6144[4742] = cin[4906];
assign cj_6144[4743] = cin[5265];
assign cj_6144[4744] = cin[440];
assign cj_6144[4745] = cin[2719];
assign cj_6144[4746] = cin[5958];
assign cj_6144[4747] = cin[4013];
assign cj_6144[4748] = cin[3028];
assign cj_6144[4749] = cin[3003];
assign cj_6144[4750] = cin[3938];
assign cj_6144[4751] = cin[5833];
assign cj_6144[4752] = cin[2544];
assign cj_6144[4753] = cin[215];
assign cj_6144[4754] = cin[4990];
assign cj_6144[4755] = cin[4581];
assign cj_6144[4756] = cin[5132];
assign cj_6144[4757] = cin[499];
assign cj_6144[4758] = cin[2970];
assign cj_6144[4759] = cin[257];
assign cj_6144[4760] = cin[4648];
assign cj_6144[4761] = cin[3855];
assign cj_6144[4762] = cin[4022];
assign cj_6144[4763] = cin[5149];
assign cj_6144[4764] = cin[1092];
assign cj_6144[4765] = cin[4139];
assign cj_6144[4766] = cin[2002];
assign cj_6144[4767] = cin[825];
assign cj_6144[4768] = cin[608];
assign cj_6144[4769] = cin[1351];
assign cj_6144[4770] = cin[3054];
assign cj_6144[4771] = cin[5717];
assign cj_6144[4772] = cin[3196];
assign cj_6144[4773] = cin[1635];
assign cj_6144[4774] = cin[1034];
assign cj_6144[4775] = cin[1393];
assign cj_6144[4776] = cin[2712];
assign cj_6144[4777] = cin[4991];
assign cj_6144[4778] = cin[2086];
assign cj_6144[4779] = cin[141];
assign cj_6144[4780] = cin[5300];
assign cj_6144[4781] = cin[5275];
assign cj_6144[4782] = cin[66];
assign cj_6144[4783] = cin[1961];
assign cj_6144[4784] = cin[4816];
assign cj_6144[4785] = cin[2487];
assign cj_6144[4786] = cin[1118];
assign cj_6144[4787] = cin[709];
assign cj_6144[4788] = cin[1260];
assign cj_6144[4789] = cin[2771];
assign cj_6144[4790] = cin[5242];
assign cj_6144[4791] = cin[2529];
assign cj_6144[4792] = cin[776];
assign cj_6144[4793] = cin[6127];
assign cj_6144[4794] = cin[150];
assign cj_6144[4795] = cin[1277];
assign cj_6144[4796] = cin[3364];
assign cj_6144[4797] = cin[267];
assign cj_6144[4798] = cin[4274];
assign cj_6144[4799] = cin[3097];
assign cj_6144[4800] = cin[2880];
assign cj_6144[4801] = cin[3623];
assign cj_6144[4802] = cin[5326];
assign cj_6144[4803] = cin[1845];
assign cj_6144[4804] = cin[5468];
assign cj_6144[4805] = cin[3907];
assign cj_6144[4806] = cin[3306];
assign cj_6144[4807] = cin[3665];
assign cj_6144[4808] = cin[4984];
assign cj_6144[4809] = cin[1119];
assign cj_6144[4810] = cin[4358];
assign cj_6144[4811] = cin[2413];
assign cj_6144[4812] = cin[1428];
assign cj_6144[4813] = cin[1403];
assign cj_6144[4814] = cin[2338];
assign cj_6144[4815] = cin[4233];
assign cj_6144[4816] = cin[944];
assign cj_6144[4817] = cin[4759];
assign cj_6144[4818] = cin[3390];
assign cj_6144[4819] = cin[2981];
assign cj_6144[4820] = cin[3532];
assign cj_6144[4821] = cin[5043];
assign cj_6144[4822] = cin[1370];
assign cj_6144[4823] = cin[4801];
assign cj_6144[4824] = cin[3048];
assign cj_6144[4825] = cin[2255];
assign cj_6144[4826] = cin[2422];
assign cj_6144[4827] = cin[3549];
assign cj_6144[4828] = cin[5636];
assign cj_6144[4829] = cin[2539];
assign cj_6144[4830] = cin[402];
assign cj_6144[4831] = cin[5369];
assign cj_6144[4832] = cin[5152];
assign cj_6144[4833] = cin[5895];
assign cj_6144[4834] = cin[1454];
assign cj_6144[4835] = cin[4117];
assign cj_6144[4836] = cin[1596];
assign cj_6144[4837] = cin[35];
assign cj_6144[4838] = cin[5578];
assign cj_6144[4839] = cin[5937];
assign cj_6144[4840] = cin[1112];
assign cj_6144[4841] = cin[3391];
assign cj_6144[4842] = cin[486];
assign cj_6144[4843] = cin[4685];
assign cj_6144[4844] = cin[3700];
assign cj_6144[4845] = cin[3675];
assign cj_6144[4846] = cin[4610];
assign cj_6144[4847] = cin[361];
assign cj_6144[4848] = cin[3216];
assign cj_6144[4849] = cin[887];
assign cj_6144[4850] = cin[5662];
assign cj_6144[4851] = cin[5253];
assign cj_6144[4852] = cin[5804];
assign cj_6144[4853] = cin[1171];
assign cj_6144[4854] = cin[3642];
assign cj_6144[4855] = cin[929];
assign cj_6144[4856] = cin[5320];
assign cj_6144[4857] = cin[4527];
assign cj_6144[4858] = cin[4694];
assign cj_6144[4859] = cin[5821];
assign cj_6144[4860] = cin[1764];
assign cj_6144[4861] = cin[4811];
assign cj_6144[4862] = cin[2674];
assign cj_6144[4863] = cin[1497];
assign cj_6144[4864] = cin[1280];
assign cj_6144[4865] = cin[2023];
assign cj_6144[4866] = cin[3726];
assign cj_6144[4867] = cin[245];
assign cj_6144[4868] = cin[3868];
assign cj_6144[4869] = cin[2307];
assign cj_6144[4870] = cin[1706];
assign cj_6144[4871] = cin[2065];
assign cj_6144[4872] = cin[3384];
assign cj_6144[4873] = cin[5663];
assign cj_6144[4874] = cin[2758];
assign cj_6144[4875] = cin[813];
assign cj_6144[4876] = cin[5972];
assign cj_6144[4877] = cin[5947];
assign cj_6144[4878] = cin[738];
assign cj_6144[4879] = cin[2633];
assign cj_6144[4880] = cin[5488];
assign cj_6144[4881] = cin[3159];
assign cj_6144[4882] = cin[1790];
assign cj_6144[4883] = cin[1381];
assign cj_6144[4884] = cin[1932];
assign cj_6144[4885] = cin[3443];
assign cj_6144[4886] = cin[5914];
assign cj_6144[4887] = cin[3201];
assign cj_6144[4888] = cin[1448];
assign cj_6144[4889] = cin[655];
assign cj_6144[4890] = cin[822];
assign cj_6144[4891] = cin[1949];
assign cj_6144[4892] = cin[4036];
assign cj_6144[4893] = cin[939];
assign cj_6144[4894] = cin[4946];
assign cj_6144[4895] = cin[3769];
assign cj_6144[4896] = cin[3552];
assign cj_6144[4897] = cin[4295];
assign cj_6144[4898] = cin[5998];
assign cj_6144[4899] = cin[2517];
assign cj_6144[4900] = cin[6140];
assign cj_6144[4901] = cin[4579];
assign cj_6144[4902] = cin[3978];
assign cj_6144[4903] = cin[4337];
assign cj_6144[4904] = cin[5656];
assign cj_6144[4905] = cin[1791];
assign cj_6144[4906] = cin[5030];
assign cj_6144[4907] = cin[3085];
assign cj_6144[4908] = cin[2100];
assign cj_6144[4909] = cin[2075];
assign cj_6144[4910] = cin[3010];
assign cj_6144[4911] = cin[4905];
assign cj_6144[4912] = cin[1616];
assign cj_6144[4913] = cin[5431];
assign cj_6144[4914] = cin[4062];
assign cj_6144[4915] = cin[3653];
assign cj_6144[4916] = cin[4204];
assign cj_6144[4917] = cin[5715];
assign cj_6144[4918] = cin[2042];
assign cj_6144[4919] = cin[5473];
assign cj_6144[4920] = cin[3720];
assign cj_6144[4921] = cin[2927];
assign cj_6144[4922] = cin[3094];
assign cj_6144[4923] = cin[4221];
assign cj_6144[4924] = cin[164];
assign cj_6144[4925] = cin[3211];
assign cj_6144[4926] = cin[1074];
assign cj_6144[4927] = cin[6041];
assign cj_6144[4928] = cin[5824];
assign cj_6144[4929] = cin[423];
assign cj_6144[4930] = cin[2126];
assign cj_6144[4931] = cin[4789];
assign cj_6144[4932] = cin[2268];
assign cj_6144[4933] = cin[707];
assign cj_6144[4934] = cin[106];
assign cj_6144[4935] = cin[465];
assign cj_6144[4936] = cin[1784];
assign cj_6144[4937] = cin[4063];
assign cj_6144[4938] = cin[1158];
assign cj_6144[4939] = cin[5357];
assign cj_6144[4940] = cin[4372];
assign cj_6144[4941] = cin[4347];
assign cj_6144[4942] = cin[5282];
assign cj_6144[4943] = cin[1033];
assign cj_6144[4944] = cin[3888];
assign cj_6144[4945] = cin[1559];
assign cj_6144[4946] = cin[190];
assign cj_6144[4947] = cin[5925];
assign cj_6144[4948] = cin[332];
assign cj_6144[4949] = cin[1843];
assign cj_6144[4950] = cin[4314];
assign cj_6144[4951] = cin[1601];
assign cj_6144[4952] = cin[5992];
assign cj_6144[4953] = cin[5199];
assign cj_6144[4954] = cin[5366];
assign cj_6144[4955] = cin[349];
assign cj_6144[4956] = cin[2436];
assign cj_6144[4957] = cin[5483];
assign cj_6144[4958] = cin[3346];
assign cj_6144[4959] = cin[2169];
assign cj_6144[4960] = cin[1952];
assign cj_6144[4961] = cin[2695];
assign cj_6144[4962] = cin[4398];
assign cj_6144[4963] = cin[917];
assign cj_6144[4964] = cin[4540];
assign cj_6144[4965] = cin[2979];
assign cj_6144[4966] = cin[2378];
assign cj_6144[4967] = cin[2737];
assign cj_6144[4968] = cin[4056];
assign cj_6144[4969] = cin[191];
assign cj_6144[4970] = cin[3430];
assign cj_6144[4971] = cin[1485];
assign cj_6144[4972] = cin[500];
assign cj_6144[4973] = cin[475];
assign cj_6144[4974] = cin[1410];
assign cj_6144[4975] = cin[3305];
assign cj_6144[4976] = cin[16];
assign cj_6144[4977] = cin[3831];
assign cj_6144[4978] = cin[2462];
assign cj_6144[4979] = cin[2053];
assign cj_6144[4980] = cin[2604];
assign cj_6144[4981] = cin[4115];
assign cj_6144[4982] = cin[442];
assign cj_6144[4983] = cin[3873];
assign cj_6144[4984] = cin[2120];
assign cj_6144[4985] = cin[1327];
assign cj_6144[4986] = cin[1494];
assign cj_6144[4987] = cin[2621];
assign cj_6144[4988] = cin[4708];
assign cj_6144[4989] = cin[1611];
assign cj_6144[4990] = cin[5618];
assign cj_6144[4991] = cin[4441];
assign cj_6144[4992] = cin[4224];
assign cj_6144[4993] = cin[4967];
assign cj_6144[4994] = cin[526];
assign cj_6144[4995] = cin[3189];
assign cj_6144[4996] = cin[668];
assign cj_6144[4997] = cin[5251];
assign cj_6144[4998] = cin[4650];
assign cj_6144[4999] = cin[5009];
assign cj_6144[5000] = cin[184];
assign cj_6144[5001] = cin[2463];
assign cj_6144[5002] = cin[5702];
assign cj_6144[5003] = cin[3757];
assign cj_6144[5004] = cin[2772];
assign cj_6144[5005] = cin[2747];
assign cj_6144[5006] = cin[3682];
assign cj_6144[5007] = cin[5577];
assign cj_6144[5008] = cin[2288];
assign cj_6144[5009] = cin[6103];
assign cj_6144[5010] = cin[4734];
assign cj_6144[5011] = cin[4325];
assign cj_6144[5012] = cin[4876];
assign cj_6144[5013] = cin[243];
assign cj_6144[5014] = cin[2714];
assign cj_6144[5015] = cin[1];
assign cj_6144[5016] = cin[4392];
assign cj_6144[5017] = cin[3599];
assign cj_6144[5018] = cin[3766];
assign cj_6144[5019] = cin[4893];
assign cj_6144[5020] = cin[836];
assign cj_6144[5021] = cin[3883];
assign cj_6144[5022] = cin[1746];
assign cj_6144[5023] = cin[569];
assign cj_6144[5024] = cin[352];
assign cj_6144[5025] = cin[1095];
assign cj_6144[5026] = cin[2798];
assign cj_6144[5027] = cin[5461];
assign cj_6144[5028] = cin[2940];
assign cj_6144[5029] = cin[1379];
assign cj_6144[5030] = cin[778];
assign cj_6144[5031] = cin[1137];
assign cj_6144[5032] = cin[2456];
assign cj_6144[5033] = cin[4735];
assign cj_6144[5034] = cin[1830];
assign cj_6144[5035] = cin[6029];
assign cj_6144[5036] = cin[5044];
assign cj_6144[5037] = cin[5019];
assign cj_6144[5038] = cin[5954];
assign cj_6144[5039] = cin[1705];
assign cj_6144[5040] = cin[4560];
assign cj_6144[5041] = cin[2231];
assign cj_6144[5042] = cin[862];
assign cj_6144[5043] = cin[453];
assign cj_6144[5044] = cin[1004];
assign cj_6144[5045] = cin[2515];
assign cj_6144[5046] = cin[4986];
assign cj_6144[5047] = cin[2273];
assign cj_6144[5048] = cin[520];
assign cj_6144[5049] = cin[5871];
assign cj_6144[5050] = cin[6038];
assign cj_6144[5051] = cin[1021];
assign cj_6144[5052] = cin[3108];
assign cj_6144[5053] = cin[11];
assign cj_6144[5054] = cin[4018];
assign cj_6144[5055] = cin[2841];
assign cj_6144[5056] = cin[2624];
assign cj_6144[5057] = cin[3367];
assign cj_6144[5058] = cin[5070];
assign cj_6144[5059] = cin[1589];
assign cj_6144[5060] = cin[5212];
assign cj_6144[5061] = cin[3651];
assign cj_6144[5062] = cin[3050];
assign cj_6144[5063] = cin[3409];
assign cj_6144[5064] = cin[4728];
assign cj_6144[5065] = cin[863];
assign cj_6144[5066] = cin[4102];
assign cj_6144[5067] = cin[2157];
assign cj_6144[5068] = cin[1172];
assign cj_6144[5069] = cin[1147];
assign cj_6144[5070] = cin[2082];
assign cj_6144[5071] = cin[3977];
assign cj_6144[5072] = cin[688];
assign cj_6144[5073] = cin[4503];
assign cj_6144[5074] = cin[3134];
assign cj_6144[5075] = cin[2725];
assign cj_6144[5076] = cin[3276];
assign cj_6144[5077] = cin[4787];
assign cj_6144[5078] = cin[1114];
assign cj_6144[5079] = cin[4545];
assign cj_6144[5080] = cin[2792];
assign cj_6144[5081] = cin[1999];
assign cj_6144[5082] = cin[2166];
assign cj_6144[5083] = cin[3293];
assign cj_6144[5084] = cin[5380];
assign cj_6144[5085] = cin[2283];
assign cj_6144[5086] = cin[146];
assign cj_6144[5087] = cin[5113];
assign cj_6144[5088] = cin[4896];
assign cj_6144[5089] = cin[5639];
assign cj_6144[5090] = cin[1198];
assign cj_6144[5091] = cin[3861];
assign cj_6144[5092] = cin[1340];
assign cj_6144[5093] = cin[5923];
assign cj_6144[5094] = cin[5322];
assign cj_6144[5095] = cin[5681];
assign cj_6144[5096] = cin[856];
assign cj_6144[5097] = cin[3135];
assign cj_6144[5098] = cin[230];
assign cj_6144[5099] = cin[4429];
assign cj_6144[5100] = cin[3444];
assign cj_6144[5101] = cin[3419];
assign cj_6144[5102] = cin[4354];
assign cj_6144[5103] = cin[105];
assign cj_6144[5104] = cin[2960];
assign cj_6144[5105] = cin[631];
assign cj_6144[5106] = cin[5406];
assign cj_6144[5107] = cin[4997];
assign cj_6144[5108] = cin[5548];
assign cj_6144[5109] = cin[915];
assign cj_6144[5110] = cin[3386];
assign cj_6144[5111] = cin[673];
assign cj_6144[5112] = cin[5064];
assign cj_6144[5113] = cin[4271];
assign cj_6144[5114] = cin[4438];
assign cj_6144[5115] = cin[5565];
assign cj_6144[5116] = cin[1508];
assign cj_6144[5117] = cin[4555];
assign cj_6144[5118] = cin[2418];
assign cj_6144[5119] = cin[1241];
assign cj_6144[5120] = cin[1024];
assign cj_6144[5121] = cin[1767];
assign cj_6144[5122] = cin[3470];
assign cj_6144[5123] = cin[6133];
assign cj_6144[5124] = cin[3612];
assign cj_6144[5125] = cin[2051];
assign cj_6144[5126] = cin[1450];
assign cj_6144[5127] = cin[1809];
assign cj_6144[5128] = cin[3128];
assign cj_6144[5129] = cin[5407];
assign cj_6144[5130] = cin[2502];
assign cj_6144[5131] = cin[557];
assign cj_6144[5132] = cin[5716];
assign cj_6144[5133] = cin[5691];
assign cj_6144[5134] = cin[482];
assign cj_6144[5135] = cin[2377];
assign cj_6144[5136] = cin[5232];
assign cj_6144[5137] = cin[2903];
assign cj_6144[5138] = cin[1534];
assign cj_6144[5139] = cin[1125];
assign cj_6144[5140] = cin[1676];
assign cj_6144[5141] = cin[3187];
assign cj_6144[5142] = cin[5658];
assign cj_6144[5143] = cin[2945];
assign cj_6144[5144] = cin[1192];
assign cj_6144[5145] = cin[399];
assign cj_6144[5146] = cin[566];
assign cj_6144[5147] = cin[1693];
assign cj_6144[5148] = cin[3780];
assign cj_6144[5149] = cin[683];
assign cj_6144[5150] = cin[4690];
assign cj_6144[5151] = cin[3513];
assign cj_6144[5152] = cin[3296];
assign cj_6144[5153] = cin[4039];
assign cj_6144[5154] = cin[5742];
assign cj_6144[5155] = cin[2261];
assign cj_6144[5156] = cin[5884];
assign cj_6144[5157] = cin[4323];
assign cj_6144[5158] = cin[3722];
assign cj_6144[5159] = cin[4081];
assign cj_6144[5160] = cin[5400];
assign cj_6144[5161] = cin[1535];
assign cj_6144[5162] = cin[4774];
assign cj_6144[5163] = cin[2829];
assign cj_6144[5164] = cin[1844];
assign cj_6144[5165] = cin[1819];
assign cj_6144[5166] = cin[2754];
assign cj_6144[5167] = cin[4649];
assign cj_6144[5168] = cin[1360];
assign cj_6144[5169] = cin[5175];
assign cj_6144[5170] = cin[3806];
assign cj_6144[5171] = cin[3397];
assign cj_6144[5172] = cin[3948];
assign cj_6144[5173] = cin[5459];
assign cj_6144[5174] = cin[1786];
assign cj_6144[5175] = cin[5217];
assign cj_6144[5176] = cin[3464];
assign cj_6144[5177] = cin[2671];
assign cj_6144[5178] = cin[2838];
assign cj_6144[5179] = cin[3965];
assign cj_6144[5180] = cin[6052];
assign cj_6144[5181] = cin[2955];
assign cj_6144[5182] = cin[818];
assign cj_6144[5183] = cin[5785];
assign cj_6144[5184] = cin[5568];
assign cj_6144[5185] = cin[167];
assign cj_6144[5186] = cin[1870];
assign cj_6144[5187] = cin[4533];
assign cj_6144[5188] = cin[2012];
assign cj_6144[5189] = cin[451];
assign cj_6144[5190] = cin[5994];
assign cj_6144[5191] = cin[209];
assign cj_6144[5192] = cin[1528];
assign cj_6144[5193] = cin[3807];
assign cj_6144[5194] = cin[902];
assign cj_6144[5195] = cin[5101];
assign cj_6144[5196] = cin[4116];
assign cj_6144[5197] = cin[4091];
assign cj_6144[5198] = cin[5026];
assign cj_6144[5199] = cin[777];
assign cj_6144[5200] = cin[3632];
assign cj_6144[5201] = cin[1303];
assign cj_6144[5202] = cin[6078];
assign cj_6144[5203] = cin[5669];
assign cj_6144[5204] = cin[76];
assign cj_6144[5205] = cin[1587];
assign cj_6144[5206] = cin[4058];
assign cj_6144[5207] = cin[1345];
assign cj_6144[5208] = cin[5736];
assign cj_6144[5209] = cin[4943];
assign cj_6144[5210] = cin[5110];
assign cj_6144[5211] = cin[93];
assign cj_6144[5212] = cin[2180];
assign cj_6144[5213] = cin[5227];
assign cj_6144[5214] = cin[3090];
assign cj_6144[5215] = cin[1913];
assign cj_6144[5216] = cin[1696];
assign cj_6144[5217] = cin[2439];
assign cj_6144[5218] = cin[4142];
assign cj_6144[5219] = cin[661];
assign cj_6144[5220] = cin[4284];
assign cj_6144[5221] = cin[2723];
assign cj_6144[5222] = cin[2122];
assign cj_6144[5223] = cin[2481];
assign cj_6144[5224] = cin[3800];
assign cj_6144[5225] = cin[6079];
assign cj_6144[5226] = cin[3174];
assign cj_6144[5227] = cin[1229];
assign cj_6144[5228] = cin[244];
assign cj_6144[5229] = cin[219];
assign cj_6144[5230] = cin[1154];
assign cj_6144[5231] = cin[3049];
assign cj_6144[5232] = cin[5904];
assign cj_6144[5233] = cin[3575];
assign cj_6144[5234] = cin[2206];
assign cj_6144[5235] = cin[1797];
assign cj_6144[5236] = cin[2348];
assign cj_6144[5237] = cin[3859];
assign cj_6144[5238] = cin[186];
assign cj_6144[5239] = cin[3617];
assign cj_6144[5240] = cin[1864];
assign cj_6144[5241] = cin[1071];
assign cj_6144[5242] = cin[1238];
assign cj_6144[5243] = cin[2365];
assign cj_6144[5244] = cin[4452];
assign cj_6144[5245] = cin[1355];
assign cj_6144[5246] = cin[5362];
assign cj_6144[5247] = cin[4185];
assign cj_6144[5248] = cin[3968];
assign cj_6144[5249] = cin[4711];
assign cj_6144[5250] = cin[270];
assign cj_6144[5251] = cin[2933];
assign cj_6144[5252] = cin[412];
assign cj_6144[5253] = cin[4995];
assign cj_6144[5254] = cin[4394];
assign cj_6144[5255] = cin[4753];
assign cj_6144[5256] = cin[6072];
assign cj_6144[5257] = cin[2207];
assign cj_6144[5258] = cin[5446];
assign cj_6144[5259] = cin[3501];
assign cj_6144[5260] = cin[2516];
assign cj_6144[5261] = cin[2491];
assign cj_6144[5262] = cin[3426];
assign cj_6144[5263] = cin[5321];
assign cj_6144[5264] = cin[2032];
assign cj_6144[5265] = cin[5847];
assign cj_6144[5266] = cin[4478];
assign cj_6144[5267] = cin[4069];
assign cj_6144[5268] = cin[4620];
assign cj_6144[5269] = cin[6131];
assign cj_6144[5270] = cin[2458];
assign cj_6144[5271] = cin[5889];
assign cj_6144[5272] = cin[4136];
assign cj_6144[5273] = cin[3343];
assign cj_6144[5274] = cin[3510];
assign cj_6144[5275] = cin[4637];
assign cj_6144[5276] = cin[580];
assign cj_6144[5277] = cin[3627];
assign cj_6144[5278] = cin[1490];
assign cj_6144[5279] = cin[313];
assign cj_6144[5280] = cin[96];
assign cj_6144[5281] = cin[839];
assign cj_6144[5282] = cin[2542];
assign cj_6144[5283] = cin[5205];
assign cj_6144[5284] = cin[2684];
assign cj_6144[5285] = cin[1123];
assign cj_6144[5286] = cin[522];
assign cj_6144[5287] = cin[881];
assign cj_6144[5288] = cin[2200];
assign cj_6144[5289] = cin[4479];
assign cj_6144[5290] = cin[1574];
assign cj_6144[5291] = cin[5773];
assign cj_6144[5292] = cin[4788];
assign cj_6144[5293] = cin[4763];
assign cj_6144[5294] = cin[5698];
assign cj_6144[5295] = cin[1449];
assign cj_6144[5296] = cin[4304];
assign cj_6144[5297] = cin[1975];
assign cj_6144[5298] = cin[606];
assign cj_6144[5299] = cin[197];
assign cj_6144[5300] = cin[748];
assign cj_6144[5301] = cin[2259];
assign cj_6144[5302] = cin[4730];
assign cj_6144[5303] = cin[2017];
assign cj_6144[5304] = cin[264];
assign cj_6144[5305] = cin[5615];
assign cj_6144[5306] = cin[5782];
assign cj_6144[5307] = cin[765];
assign cj_6144[5308] = cin[2852];
assign cj_6144[5309] = cin[5899];
assign cj_6144[5310] = cin[3762];
assign cj_6144[5311] = cin[2585];
assign cj_6144[5312] = cin[2368];
assign cj_6144[5313] = cin[3111];
assign cj_6144[5314] = cin[4814];
assign cj_6144[5315] = cin[1333];
assign cj_6144[5316] = cin[4956];
assign cj_6144[5317] = cin[3395];
assign cj_6144[5318] = cin[2794];
assign cj_6144[5319] = cin[3153];
assign cj_6144[5320] = cin[4472];
assign cj_6144[5321] = cin[607];
assign cj_6144[5322] = cin[3846];
assign cj_6144[5323] = cin[1901];
assign cj_6144[5324] = cin[916];
assign cj_6144[5325] = cin[891];
assign cj_6144[5326] = cin[1826];
assign cj_6144[5327] = cin[3721];
assign cj_6144[5328] = cin[432];
assign cj_6144[5329] = cin[4247];
assign cj_6144[5330] = cin[2878];
assign cj_6144[5331] = cin[2469];
assign cj_6144[5332] = cin[3020];
assign cj_6144[5333] = cin[4531];
assign cj_6144[5334] = cin[858];
assign cj_6144[5335] = cin[4289];
assign cj_6144[5336] = cin[2536];
assign cj_6144[5337] = cin[1743];
assign cj_6144[5338] = cin[1910];
assign cj_6144[5339] = cin[3037];
assign cj_6144[5340] = cin[5124];
assign cj_6144[5341] = cin[2027];
assign cj_6144[5342] = cin[6034];
assign cj_6144[5343] = cin[4857];
assign cj_6144[5344] = cin[4640];
assign cj_6144[5345] = cin[5383];
assign cj_6144[5346] = cin[942];
assign cj_6144[5347] = cin[3605];
assign cj_6144[5348] = cin[1084];
assign cj_6144[5349] = cin[5667];
assign cj_6144[5350] = cin[5066];
assign cj_6144[5351] = cin[5425];
assign cj_6144[5352] = cin[600];
assign cj_6144[5353] = cin[2879];
assign cj_6144[5354] = cin[6118];
assign cj_6144[5355] = cin[4173];
assign cj_6144[5356] = cin[3188];
assign cj_6144[5357] = cin[3163];
assign cj_6144[5358] = cin[4098];
assign cj_6144[5359] = cin[5993];
assign cj_6144[5360] = cin[2704];
assign cj_6144[5361] = cin[375];
assign cj_6144[5362] = cin[5150];
assign cj_6144[5363] = cin[4741];
assign cj_6144[5364] = cin[5292];
assign cj_6144[5365] = cin[659];
assign cj_6144[5366] = cin[3130];
assign cj_6144[5367] = cin[417];
assign cj_6144[5368] = cin[4808];
assign cj_6144[5369] = cin[4015];
assign cj_6144[5370] = cin[4182];
assign cj_6144[5371] = cin[5309];
assign cj_6144[5372] = cin[1252];
assign cj_6144[5373] = cin[4299];
assign cj_6144[5374] = cin[2162];
assign cj_6144[5375] = cin[985];
assign cj_6144[5376] = cin[768];
assign cj_6144[5377] = cin[1511];
assign cj_6144[5378] = cin[3214];
assign cj_6144[5379] = cin[5877];
assign cj_6144[5380] = cin[3356];
assign cj_6144[5381] = cin[1795];
assign cj_6144[5382] = cin[1194];
assign cj_6144[5383] = cin[1553];
assign cj_6144[5384] = cin[2872];
assign cj_6144[5385] = cin[5151];
assign cj_6144[5386] = cin[2246];
assign cj_6144[5387] = cin[301];
assign cj_6144[5388] = cin[5460];
assign cj_6144[5389] = cin[5435];
assign cj_6144[5390] = cin[226];
assign cj_6144[5391] = cin[2121];
assign cj_6144[5392] = cin[4976];
assign cj_6144[5393] = cin[2647];
assign cj_6144[5394] = cin[1278];
assign cj_6144[5395] = cin[869];
assign cj_6144[5396] = cin[1420];
assign cj_6144[5397] = cin[2931];
assign cj_6144[5398] = cin[5402];
assign cj_6144[5399] = cin[2689];
assign cj_6144[5400] = cin[936];
assign cj_6144[5401] = cin[143];
assign cj_6144[5402] = cin[310];
assign cj_6144[5403] = cin[1437];
assign cj_6144[5404] = cin[3524];
assign cj_6144[5405] = cin[427];
assign cj_6144[5406] = cin[4434];
assign cj_6144[5407] = cin[3257];
assign cj_6144[5408] = cin[3040];
assign cj_6144[5409] = cin[3783];
assign cj_6144[5410] = cin[5486];
assign cj_6144[5411] = cin[2005];
assign cj_6144[5412] = cin[5628];
assign cj_6144[5413] = cin[4067];
assign cj_6144[5414] = cin[3466];
assign cj_6144[5415] = cin[3825];
assign cj_6144[5416] = cin[5144];
assign cj_6144[5417] = cin[1279];
assign cj_6144[5418] = cin[4518];
assign cj_6144[5419] = cin[2573];
assign cj_6144[5420] = cin[1588];
assign cj_6144[5421] = cin[1563];
assign cj_6144[5422] = cin[2498];
assign cj_6144[5423] = cin[4393];
assign cj_6144[5424] = cin[1104];
assign cj_6144[5425] = cin[4919];
assign cj_6144[5426] = cin[3550];
assign cj_6144[5427] = cin[3141];
assign cj_6144[5428] = cin[3692];
assign cj_6144[5429] = cin[5203];
assign cj_6144[5430] = cin[1530];
assign cj_6144[5431] = cin[4961];
assign cj_6144[5432] = cin[3208];
assign cj_6144[5433] = cin[2415];
assign cj_6144[5434] = cin[2582];
assign cj_6144[5435] = cin[3709];
assign cj_6144[5436] = cin[5796];
assign cj_6144[5437] = cin[2699];
assign cj_6144[5438] = cin[562];
assign cj_6144[5439] = cin[5529];
assign cj_6144[5440] = cin[5312];
assign cj_6144[5441] = cin[6055];
assign cj_6144[5442] = cin[1614];
assign cj_6144[5443] = cin[4277];
assign cj_6144[5444] = cin[1756];
assign cj_6144[5445] = cin[195];
assign cj_6144[5446] = cin[5738];
assign cj_6144[5447] = cin[6097];
assign cj_6144[5448] = cin[1272];
assign cj_6144[5449] = cin[3551];
assign cj_6144[5450] = cin[646];
assign cj_6144[5451] = cin[4845];
assign cj_6144[5452] = cin[3860];
assign cj_6144[5453] = cin[3835];
assign cj_6144[5454] = cin[4770];
assign cj_6144[5455] = cin[521];
assign cj_6144[5456] = cin[3376];
assign cj_6144[5457] = cin[1047];
assign cj_6144[5458] = cin[5822];
assign cj_6144[5459] = cin[5413];
assign cj_6144[5460] = cin[5964];
assign cj_6144[5461] = cin[1331];
assign cj_6144[5462] = cin[3802];
assign cj_6144[5463] = cin[1089];
assign cj_6144[5464] = cin[5480];
assign cj_6144[5465] = cin[4687];
assign cj_6144[5466] = cin[4854];
assign cj_6144[5467] = cin[5981];
assign cj_6144[5468] = cin[1924];
assign cj_6144[5469] = cin[4971];
assign cj_6144[5470] = cin[2834];
assign cj_6144[5471] = cin[1657];
assign cj_6144[5472] = cin[1440];
assign cj_6144[5473] = cin[2183];
assign cj_6144[5474] = cin[3886];
assign cj_6144[5475] = cin[405];
assign cj_6144[5476] = cin[4028];
assign cj_6144[5477] = cin[2467];
assign cj_6144[5478] = cin[1866];
assign cj_6144[5479] = cin[2225];
assign cj_6144[5480] = cin[3544];
assign cj_6144[5481] = cin[5823];
assign cj_6144[5482] = cin[2918];
assign cj_6144[5483] = cin[973];
assign cj_6144[5484] = cin[6132];
assign cj_6144[5485] = cin[6107];
assign cj_6144[5486] = cin[898];
assign cj_6144[5487] = cin[2793];
assign cj_6144[5488] = cin[5648];
assign cj_6144[5489] = cin[3319];
assign cj_6144[5490] = cin[1950];
assign cj_6144[5491] = cin[1541];
assign cj_6144[5492] = cin[2092];
assign cj_6144[5493] = cin[3603];
assign cj_6144[5494] = cin[6074];
assign cj_6144[5495] = cin[3361];
assign cj_6144[5496] = cin[1608];
assign cj_6144[5497] = cin[815];
assign cj_6144[5498] = cin[982];
assign cj_6144[5499] = cin[2109];
assign cj_6144[5500] = cin[4196];
assign cj_6144[5501] = cin[1099];
assign cj_6144[5502] = cin[5106];
assign cj_6144[5503] = cin[3929];
assign cj_6144[5504] = cin[3712];
assign cj_6144[5505] = cin[4455];
assign cj_6144[5506] = cin[14];
assign cj_6144[5507] = cin[2677];
assign cj_6144[5508] = cin[156];
assign cj_6144[5509] = cin[4739];
assign cj_6144[5510] = cin[4138];
assign cj_6144[5511] = cin[4497];
assign cj_6144[5512] = cin[5816];
assign cj_6144[5513] = cin[1951];
assign cj_6144[5514] = cin[5190];
assign cj_6144[5515] = cin[3245];
assign cj_6144[5516] = cin[2260];
assign cj_6144[5517] = cin[2235];
assign cj_6144[5518] = cin[3170];
assign cj_6144[5519] = cin[5065];
assign cj_6144[5520] = cin[1776];
assign cj_6144[5521] = cin[5591];
assign cj_6144[5522] = cin[4222];
assign cj_6144[5523] = cin[3813];
assign cj_6144[5524] = cin[4364];
assign cj_6144[5525] = cin[5875];
assign cj_6144[5526] = cin[2202];
assign cj_6144[5527] = cin[5633];
assign cj_6144[5528] = cin[3880];
assign cj_6144[5529] = cin[3087];
assign cj_6144[5530] = cin[3254];
assign cj_6144[5531] = cin[4381];
assign cj_6144[5532] = cin[324];
assign cj_6144[5533] = cin[3371];
assign cj_6144[5534] = cin[1234];
assign cj_6144[5535] = cin[57];
assign cj_6144[5536] = cin[5984];
assign cj_6144[5537] = cin[583];
assign cj_6144[5538] = cin[2286];
assign cj_6144[5539] = cin[4949];
assign cj_6144[5540] = cin[2428];
assign cj_6144[5541] = cin[867];
assign cj_6144[5542] = cin[266];
assign cj_6144[5543] = cin[625];
assign cj_6144[5544] = cin[1944];
assign cj_6144[5545] = cin[4223];
assign cj_6144[5546] = cin[1318];
assign cj_6144[5547] = cin[5517];
assign cj_6144[5548] = cin[4532];
assign cj_6144[5549] = cin[4507];
assign cj_6144[5550] = cin[5442];
assign cj_6144[5551] = cin[1193];
assign cj_6144[5552] = cin[4048];
assign cj_6144[5553] = cin[1719];
assign cj_6144[5554] = cin[350];
assign cj_6144[5555] = cin[6085];
assign cj_6144[5556] = cin[492];
assign cj_6144[5557] = cin[2003];
assign cj_6144[5558] = cin[4474];
assign cj_6144[5559] = cin[1761];
assign cj_6144[5560] = cin[8];
assign cj_6144[5561] = cin[5359];
assign cj_6144[5562] = cin[5526];
assign cj_6144[5563] = cin[509];
assign cj_6144[5564] = cin[2596];
assign cj_6144[5565] = cin[5643];
assign cj_6144[5566] = cin[3506];
assign cj_6144[5567] = cin[2329];
assign cj_6144[5568] = cin[2112];
assign cj_6144[5569] = cin[2855];
assign cj_6144[5570] = cin[4558];
assign cj_6144[5571] = cin[1077];
assign cj_6144[5572] = cin[4700];
assign cj_6144[5573] = cin[3139];
assign cj_6144[5574] = cin[2538];
assign cj_6144[5575] = cin[2897];
assign cj_6144[5576] = cin[4216];
assign cj_6144[5577] = cin[351];
assign cj_6144[5578] = cin[3590];
assign cj_6144[5579] = cin[1645];
assign cj_6144[5580] = cin[660];
assign cj_6144[5581] = cin[635];
assign cj_6144[5582] = cin[1570];
assign cj_6144[5583] = cin[3465];
assign cj_6144[5584] = cin[176];
assign cj_6144[5585] = cin[3991];
assign cj_6144[5586] = cin[2622];
assign cj_6144[5587] = cin[2213];
assign cj_6144[5588] = cin[2764];
assign cj_6144[5589] = cin[4275];
assign cj_6144[5590] = cin[602];
assign cj_6144[5591] = cin[4033];
assign cj_6144[5592] = cin[2280];
assign cj_6144[5593] = cin[1487];
assign cj_6144[5594] = cin[1654];
assign cj_6144[5595] = cin[2781];
assign cj_6144[5596] = cin[4868];
assign cj_6144[5597] = cin[1771];
assign cj_6144[5598] = cin[5778];
assign cj_6144[5599] = cin[4601];
assign cj_6144[5600] = cin[4384];
assign cj_6144[5601] = cin[5127];
assign cj_6144[5602] = cin[686];
assign cj_6144[5603] = cin[3349];
assign cj_6144[5604] = cin[828];
assign cj_6144[5605] = cin[5411];
assign cj_6144[5606] = cin[4810];
assign cj_6144[5607] = cin[5169];
assign cj_6144[5608] = cin[344];
assign cj_6144[5609] = cin[2623];
assign cj_6144[5610] = cin[5862];
assign cj_6144[5611] = cin[3917];
assign cj_6144[5612] = cin[2932];
assign cj_6144[5613] = cin[2907];
assign cj_6144[5614] = cin[3842];
assign cj_6144[5615] = cin[5737];
assign cj_6144[5616] = cin[2448];
assign cj_6144[5617] = cin[119];
assign cj_6144[5618] = cin[4894];
assign cj_6144[5619] = cin[4485];
assign cj_6144[5620] = cin[5036];
assign cj_6144[5621] = cin[403];
assign cj_6144[5622] = cin[2874];
assign cj_6144[5623] = cin[161];
assign cj_6144[5624] = cin[4552];
assign cj_6144[5625] = cin[3759];
assign cj_6144[5626] = cin[3926];
assign cj_6144[5627] = cin[5053];
assign cj_6144[5628] = cin[996];
assign cj_6144[5629] = cin[4043];
assign cj_6144[5630] = cin[1906];
assign cj_6144[5631] = cin[729];
assign cj_6144[5632] = cin[512];
assign cj_6144[5633] = cin[1255];
assign cj_6144[5634] = cin[2958];
assign cj_6144[5635] = cin[5621];
assign cj_6144[5636] = cin[3100];
assign cj_6144[5637] = cin[1539];
assign cj_6144[5638] = cin[938];
assign cj_6144[5639] = cin[1297];
assign cj_6144[5640] = cin[2616];
assign cj_6144[5641] = cin[4895];
assign cj_6144[5642] = cin[1990];
assign cj_6144[5643] = cin[45];
assign cj_6144[5644] = cin[5204];
assign cj_6144[5645] = cin[5179];
assign cj_6144[5646] = cin[6114];
assign cj_6144[5647] = cin[1865];
assign cj_6144[5648] = cin[4720];
assign cj_6144[5649] = cin[2391];
assign cj_6144[5650] = cin[1022];
assign cj_6144[5651] = cin[613];
assign cj_6144[5652] = cin[1164];
assign cj_6144[5653] = cin[2675];
assign cj_6144[5654] = cin[5146];
assign cj_6144[5655] = cin[2433];
assign cj_6144[5656] = cin[680];
assign cj_6144[5657] = cin[6031];
assign cj_6144[5658] = cin[54];
assign cj_6144[5659] = cin[1181];
assign cj_6144[5660] = cin[3268];
assign cj_6144[5661] = cin[171];
assign cj_6144[5662] = cin[4178];
assign cj_6144[5663] = cin[3001];
assign cj_6144[5664] = cin[2784];
assign cj_6144[5665] = cin[3527];
assign cj_6144[5666] = cin[5230];
assign cj_6144[5667] = cin[1749];
assign cj_6144[5668] = cin[5372];
assign cj_6144[5669] = cin[3811];
assign cj_6144[5670] = cin[3210];
assign cj_6144[5671] = cin[3569];
assign cj_6144[5672] = cin[4888];
assign cj_6144[5673] = cin[1023];
assign cj_6144[5674] = cin[4262];
assign cj_6144[5675] = cin[2317];
assign cj_6144[5676] = cin[1332];
assign cj_6144[5677] = cin[1307];
assign cj_6144[5678] = cin[2242];
assign cj_6144[5679] = cin[4137];
assign cj_6144[5680] = cin[848];
assign cj_6144[5681] = cin[4663];
assign cj_6144[5682] = cin[3294];
assign cj_6144[5683] = cin[2885];
assign cj_6144[5684] = cin[3436];
assign cj_6144[5685] = cin[4947];
assign cj_6144[5686] = cin[1274];
assign cj_6144[5687] = cin[4705];
assign cj_6144[5688] = cin[2952];
assign cj_6144[5689] = cin[2159];
assign cj_6144[5690] = cin[2326];
assign cj_6144[5691] = cin[3453];
assign cj_6144[5692] = cin[5540];
assign cj_6144[5693] = cin[2443];
assign cj_6144[5694] = cin[306];
assign cj_6144[5695] = cin[5273];
assign cj_6144[5696] = cin[5056];
assign cj_6144[5697] = cin[5799];
assign cj_6144[5698] = cin[1358];
assign cj_6144[5699] = cin[4021];
assign cj_6144[5700] = cin[1500];
assign cj_6144[5701] = cin[6083];
assign cj_6144[5702] = cin[5482];
assign cj_6144[5703] = cin[5841];
assign cj_6144[5704] = cin[1016];
assign cj_6144[5705] = cin[3295];
assign cj_6144[5706] = cin[390];
assign cj_6144[5707] = cin[4589];
assign cj_6144[5708] = cin[3604];
assign cj_6144[5709] = cin[3579];
assign cj_6144[5710] = cin[4514];
assign cj_6144[5711] = cin[265];
assign cj_6144[5712] = cin[3120];
assign cj_6144[5713] = cin[791];
assign cj_6144[5714] = cin[5566];
assign cj_6144[5715] = cin[5157];
assign cj_6144[5716] = cin[5708];
assign cj_6144[5717] = cin[1075];
assign cj_6144[5718] = cin[3546];
assign cj_6144[5719] = cin[833];
assign cj_6144[5720] = cin[5224];
assign cj_6144[5721] = cin[4431];
assign cj_6144[5722] = cin[4598];
assign cj_6144[5723] = cin[5725];
assign cj_6144[5724] = cin[1668];
assign cj_6144[5725] = cin[4715];
assign cj_6144[5726] = cin[2578];
assign cj_6144[5727] = cin[1401];
assign cj_6144[5728] = cin[1184];
assign cj_6144[5729] = cin[1927];
assign cj_6144[5730] = cin[3630];
assign cj_6144[5731] = cin[149];
assign cj_6144[5732] = cin[3772];
assign cj_6144[5733] = cin[2211];
assign cj_6144[5734] = cin[1610];
assign cj_6144[5735] = cin[1969];
assign cj_6144[5736] = cin[3288];
assign cj_6144[5737] = cin[5567];
assign cj_6144[5738] = cin[2662];
assign cj_6144[5739] = cin[717];
assign cj_6144[5740] = cin[5876];
assign cj_6144[5741] = cin[5851];
assign cj_6144[5742] = cin[642];
assign cj_6144[5743] = cin[2537];
assign cj_6144[5744] = cin[5392];
assign cj_6144[5745] = cin[3063];
assign cj_6144[5746] = cin[1694];
assign cj_6144[5747] = cin[1285];
assign cj_6144[5748] = cin[1836];
assign cj_6144[5749] = cin[3347];
assign cj_6144[5750] = cin[5818];
assign cj_6144[5751] = cin[3105];
assign cj_6144[5752] = cin[1352];
assign cj_6144[5753] = cin[559];
assign cj_6144[5754] = cin[726];
assign cj_6144[5755] = cin[1853];
assign cj_6144[5756] = cin[3940];
assign cj_6144[5757] = cin[843];
assign cj_6144[5758] = cin[4850];
assign cj_6144[5759] = cin[3673];
assign cj_6144[5760] = cin[3456];
assign cj_6144[5761] = cin[4199];
assign cj_6144[5762] = cin[5902];
assign cj_6144[5763] = cin[2421];
assign cj_6144[5764] = cin[6044];
assign cj_6144[5765] = cin[4483];
assign cj_6144[5766] = cin[3882];
assign cj_6144[5767] = cin[4241];
assign cj_6144[5768] = cin[5560];
assign cj_6144[5769] = cin[1695];
assign cj_6144[5770] = cin[4934];
assign cj_6144[5771] = cin[2989];
assign cj_6144[5772] = cin[2004];
assign cj_6144[5773] = cin[1979];
assign cj_6144[5774] = cin[2914];
assign cj_6144[5775] = cin[4809];
assign cj_6144[5776] = cin[1520];
assign cj_6144[5777] = cin[5335];
assign cj_6144[5778] = cin[3966];
assign cj_6144[5779] = cin[3557];
assign cj_6144[5780] = cin[4108];
assign cj_6144[5781] = cin[5619];
assign cj_6144[5782] = cin[1946];
assign cj_6144[5783] = cin[5377];
assign cj_6144[5784] = cin[3624];
assign cj_6144[5785] = cin[2831];
assign cj_6144[5786] = cin[2998];
assign cj_6144[5787] = cin[4125];
assign cj_6144[5788] = cin[68];
assign cj_6144[5789] = cin[3115];
assign cj_6144[5790] = cin[978];
assign cj_6144[5791] = cin[5945];
assign cj_6144[5792] = cin[5728];
assign cj_6144[5793] = cin[327];
assign cj_6144[5794] = cin[2030];
assign cj_6144[5795] = cin[4693];
assign cj_6144[5796] = cin[2172];
assign cj_6144[5797] = cin[611];
assign cj_6144[5798] = cin[10];
assign cj_6144[5799] = cin[369];
assign cj_6144[5800] = cin[1688];
assign cj_6144[5801] = cin[3967];
assign cj_6144[5802] = cin[1062];
assign cj_6144[5803] = cin[5261];
assign cj_6144[5804] = cin[4276];
assign cj_6144[5805] = cin[4251];
assign cj_6144[5806] = cin[5186];
assign cj_6144[5807] = cin[937];
assign cj_6144[5808] = cin[3792];
assign cj_6144[5809] = cin[1463];
assign cj_6144[5810] = cin[94];
assign cj_6144[5811] = cin[5829];
assign cj_6144[5812] = cin[236];
assign cj_6144[5813] = cin[1747];
assign cj_6144[5814] = cin[4218];
assign cj_6144[5815] = cin[1505];
assign cj_6144[5816] = cin[5896];
assign cj_6144[5817] = cin[5103];
assign cj_6144[5818] = cin[5270];
assign cj_6144[5819] = cin[253];
assign cj_6144[5820] = cin[2340];
assign cj_6144[5821] = cin[5387];
assign cj_6144[5822] = cin[3250];
assign cj_6144[5823] = cin[2073];
assign cj_6144[5824] = cin[1856];
assign cj_6144[5825] = cin[2599];
assign cj_6144[5826] = cin[4302];
assign cj_6144[5827] = cin[821];
assign cj_6144[5828] = cin[4444];
assign cj_6144[5829] = cin[2883];
assign cj_6144[5830] = cin[2282];
assign cj_6144[5831] = cin[2641];
assign cj_6144[5832] = cin[3960];
assign cj_6144[5833] = cin[95];
assign cj_6144[5834] = cin[3334];
assign cj_6144[5835] = cin[1389];
assign cj_6144[5836] = cin[404];
assign cj_6144[5837] = cin[379];
assign cj_6144[5838] = cin[1314];
assign cj_6144[5839] = cin[3209];
assign cj_6144[5840] = cin[6064];
assign cj_6144[5841] = cin[3735];
assign cj_6144[5842] = cin[2366];
assign cj_6144[5843] = cin[1957];
assign cj_6144[5844] = cin[2508];
assign cj_6144[5845] = cin[4019];
assign cj_6144[5846] = cin[346];
assign cj_6144[5847] = cin[3777];
assign cj_6144[5848] = cin[2024];
assign cj_6144[5849] = cin[1231];
assign cj_6144[5850] = cin[1398];
assign cj_6144[5851] = cin[2525];
assign cj_6144[5852] = cin[4612];
assign cj_6144[5853] = cin[1515];
assign cj_6144[5854] = cin[5522];
assign cj_6144[5855] = cin[4345];
assign cj_6144[5856] = cin[4128];
assign cj_6144[5857] = cin[4871];
assign cj_6144[5858] = cin[430];
assign cj_6144[5859] = cin[3093];
assign cj_6144[5860] = cin[572];
assign cj_6144[5861] = cin[5155];
assign cj_6144[5862] = cin[4554];
assign cj_6144[5863] = cin[4913];
assign cj_6144[5864] = cin[88];
assign cj_6144[5865] = cin[2367];
assign cj_6144[5866] = cin[5606];
assign cj_6144[5867] = cin[3661];
assign cj_6144[5868] = cin[2676];
assign cj_6144[5869] = cin[2651];
assign cj_6144[5870] = cin[3586];
assign cj_6144[5871] = cin[5481];
assign cj_6144[5872] = cin[2192];
assign cj_6144[5873] = cin[6007];
assign cj_6144[5874] = cin[4638];
assign cj_6144[5875] = cin[4229];
assign cj_6144[5876] = cin[4780];
assign cj_6144[5877] = cin[147];
assign cj_6144[5878] = cin[2618];
assign cj_6144[5879] = cin[6049];
assign cj_6144[5880] = cin[4296];
assign cj_6144[5881] = cin[3503];
assign cj_6144[5882] = cin[3670];
assign cj_6144[5883] = cin[4797];
assign cj_6144[5884] = cin[740];
assign cj_6144[5885] = cin[3787];
assign cj_6144[5886] = cin[1650];
assign cj_6144[5887] = cin[473];
assign cj_6144[5888] = cin[256];
assign cj_6144[5889] = cin[999];
assign cj_6144[5890] = cin[2702];
assign cj_6144[5891] = cin[5365];
assign cj_6144[5892] = cin[2844];
assign cj_6144[5893] = cin[1283];
assign cj_6144[5894] = cin[682];
assign cj_6144[5895] = cin[1041];
assign cj_6144[5896] = cin[2360];
assign cj_6144[5897] = cin[4639];
assign cj_6144[5898] = cin[1734];
assign cj_6144[5899] = cin[5933];
assign cj_6144[5900] = cin[4948];
assign cj_6144[5901] = cin[4923];
assign cj_6144[5902] = cin[5858];
assign cj_6144[5903] = cin[1609];
assign cj_6144[5904] = cin[4464];
assign cj_6144[5905] = cin[2135];
assign cj_6144[5906] = cin[766];
assign cj_6144[5907] = cin[357];
assign cj_6144[5908] = cin[908];
assign cj_6144[5909] = cin[2419];
assign cj_6144[5910] = cin[4890];
assign cj_6144[5911] = cin[2177];
assign cj_6144[5912] = cin[424];
assign cj_6144[5913] = cin[5775];
assign cj_6144[5914] = cin[5942];
assign cj_6144[5915] = cin[925];
assign cj_6144[5916] = cin[3012];
assign cj_6144[5917] = cin[6059];
assign cj_6144[5918] = cin[3922];
assign cj_6144[5919] = cin[2745];
assign cj_6144[5920] = cin[2528];
assign cj_6144[5921] = cin[3271];
assign cj_6144[5922] = cin[4974];
assign cj_6144[5923] = cin[1493];
assign cj_6144[5924] = cin[5116];
assign cj_6144[5925] = cin[3555];
assign cj_6144[5926] = cin[2954];
assign cj_6144[5927] = cin[3313];
assign cj_6144[5928] = cin[4632];
assign cj_6144[5929] = cin[767];
assign cj_6144[5930] = cin[4006];
assign cj_6144[5931] = cin[2061];
assign cj_6144[5932] = cin[1076];
assign cj_6144[5933] = cin[1051];
assign cj_6144[5934] = cin[1986];
assign cj_6144[5935] = cin[3881];
assign cj_6144[5936] = cin[592];
assign cj_6144[5937] = cin[4407];
assign cj_6144[5938] = cin[3038];
assign cj_6144[5939] = cin[2629];
assign cj_6144[5940] = cin[3180];
assign cj_6144[5941] = cin[4691];
assign cj_6144[5942] = cin[1018];
assign cj_6144[5943] = cin[4449];
assign cj_6144[5944] = cin[2696];
assign cj_6144[5945] = cin[1903];
assign cj_6144[5946] = cin[2070];
assign cj_6144[5947] = cin[3197];
assign cj_6144[5948] = cin[5284];
assign cj_6144[5949] = cin[2187];
assign cj_6144[5950] = cin[50];
assign cj_6144[5951] = cin[5017];
assign cj_6144[5952] = cin[4800];
assign cj_6144[5953] = cin[5543];
assign cj_6144[5954] = cin[1102];
assign cj_6144[5955] = cin[3765];
assign cj_6144[5956] = cin[1244];
assign cj_6144[5957] = cin[5827];
assign cj_6144[5958] = cin[5226];
assign cj_6144[5959] = cin[5585];
assign cj_6144[5960] = cin[760];
assign cj_6144[5961] = cin[3039];
assign cj_6144[5962] = cin[134];
assign cj_6144[5963] = cin[4333];
assign cj_6144[5964] = cin[3348];
assign cj_6144[5965] = cin[3323];
assign cj_6144[5966] = cin[4258];
assign cj_6144[5967] = cin[9];
assign cj_6144[5968] = cin[2864];
assign cj_6144[5969] = cin[535];
assign cj_6144[5970] = cin[5310];
assign cj_6144[5971] = cin[4901];
assign cj_6144[5972] = cin[5452];
assign cj_6144[5973] = cin[819];
assign cj_6144[5974] = cin[3290];
assign cj_6144[5975] = cin[577];
assign cj_6144[5976] = cin[4968];
assign cj_6144[5977] = cin[4175];
assign cj_6144[5978] = cin[4342];
assign cj_6144[5979] = cin[5469];
assign cj_6144[5980] = cin[1412];
assign cj_6144[5981] = cin[4459];
assign cj_6144[5982] = cin[2322];
assign cj_6144[5983] = cin[1145];
assign cj_6144[5984] = cin[928];
assign cj_6144[5985] = cin[1671];
assign cj_6144[5986] = cin[3374];
assign cj_6144[5987] = cin[6037];
assign cj_6144[5988] = cin[3516];
assign cj_6144[5989] = cin[1955];
assign cj_6144[5990] = cin[1354];
assign cj_6144[5991] = cin[1713];
assign cj_6144[5992] = cin[3032];
assign cj_6144[5993] = cin[5311];
assign cj_6144[5994] = cin[2406];
assign cj_6144[5995] = cin[461];
assign cj_6144[5996] = cin[5620];
assign cj_6144[5997] = cin[5595];
assign cj_6144[5998] = cin[386];
assign cj_6144[5999] = cin[2281];
assign cj_6144[6000] = cin[5136];
assign cj_6144[6001] = cin[2807];
assign cj_6144[6002] = cin[1438];
assign cj_6144[6003] = cin[1029];
assign cj_6144[6004] = cin[1580];
assign cj_6144[6005] = cin[3091];
assign cj_6144[6006] = cin[5562];
assign cj_6144[6007] = cin[2849];
assign cj_6144[6008] = cin[1096];
assign cj_6144[6009] = cin[303];
assign cj_6144[6010] = cin[470];
assign cj_6144[6011] = cin[1597];
assign cj_6144[6012] = cin[3684];
assign cj_6144[6013] = cin[587];
assign cj_6144[6014] = cin[4594];
assign cj_6144[6015] = cin[3417];
assign cj_6144[6016] = cin[3200];
assign cj_6144[6017] = cin[3943];
assign cj_6144[6018] = cin[5646];
assign cj_6144[6019] = cin[2165];
assign cj_6144[6020] = cin[5788];
assign cj_6144[6021] = cin[4227];
assign cj_6144[6022] = cin[3626];
assign cj_6144[6023] = cin[3985];
assign cj_6144[6024] = cin[5304];
assign cj_6144[6025] = cin[1439];
assign cj_6144[6026] = cin[4678];
assign cj_6144[6027] = cin[2733];
assign cj_6144[6028] = cin[1748];
assign cj_6144[6029] = cin[1723];
assign cj_6144[6030] = cin[2658];
assign cj_6144[6031] = cin[4553];
assign cj_6144[6032] = cin[1264];
assign cj_6144[6033] = cin[5079];
assign cj_6144[6034] = cin[3710];
assign cj_6144[6035] = cin[3301];
assign cj_6144[6036] = cin[3852];
assign cj_6144[6037] = cin[5363];
assign cj_6144[6038] = cin[1690];
assign cj_6144[6039] = cin[5121];
assign cj_6144[6040] = cin[3368];
assign cj_6144[6041] = cin[2575];
assign cj_6144[6042] = cin[2742];
assign cj_6144[6043] = cin[3869];
assign cj_6144[6044] = cin[5956];
assign cj_6144[6045] = cin[2859];
assign cj_6144[6046] = cin[722];
assign cj_6144[6047] = cin[5689];
assign cj_6144[6048] = cin[5472];
assign cj_6144[6049] = cin[71];
assign cj_6144[6050] = cin[1774];
assign cj_6144[6051] = cin[4437];
assign cj_6144[6052] = cin[1916];
assign cj_6144[6053] = cin[355];
assign cj_6144[6054] = cin[5898];
assign cj_6144[6055] = cin[113];
assign cj_6144[6056] = cin[1432];
assign cj_6144[6057] = cin[3711];
assign cj_6144[6058] = cin[806];
assign cj_6144[6059] = cin[5005];
assign cj_6144[6060] = cin[4020];
assign cj_6144[6061] = cin[3995];
assign cj_6144[6062] = cin[4930];
assign cj_6144[6063] = cin[681];
assign cj_6144[6064] = cin[3536];
assign cj_6144[6065] = cin[1207];
assign cj_6144[6066] = cin[5982];
assign cj_6144[6067] = cin[5573];
assign cj_6144[6068] = cin[6124];
assign cj_6144[6069] = cin[1491];
assign cj_6144[6070] = cin[3962];
assign cj_6144[6071] = cin[1249];
assign cj_6144[6072] = cin[5640];
assign cj_6144[6073] = cin[4847];
assign cj_6144[6074] = cin[5014];
assign cj_6144[6075] = cin[6141];
assign cj_6144[6076] = cin[2084];
assign cj_6144[6077] = cin[5131];
assign cj_6144[6078] = cin[2994];
assign cj_6144[6079] = cin[1817];
assign cj_6144[6080] = cin[1600];
assign cj_6144[6081] = cin[2343];
assign cj_6144[6082] = cin[4046];
assign cj_6144[6083] = cin[565];
assign cj_6144[6084] = cin[4188];
assign cj_6144[6085] = cin[2627];
assign cj_6144[6086] = cin[2026];
assign cj_6144[6087] = cin[2385];
assign cj_6144[6088] = cin[3704];
assign cj_6144[6089] = cin[5983];
assign cj_6144[6090] = cin[3078];
assign cj_6144[6091] = cin[1133];
assign cj_6144[6092] = cin[148];
assign cj_6144[6093] = cin[123];
assign cj_6144[6094] = cin[1058];
assign cj_6144[6095] = cin[2953];
assign cj_6144[6096] = cin[5808];
assign cj_6144[6097] = cin[3479];
assign cj_6144[6098] = cin[2110];
assign cj_6144[6099] = cin[1701];
assign cj_6144[6100] = cin[2252];
assign cj_6144[6101] = cin[3763];
assign cj_6144[6102] = cin[90];
assign cj_6144[6103] = cin[3521];
assign cj_6144[6104] = cin[1768];
assign cj_6144[6105] = cin[975];
assign cj_6144[6106] = cin[1142];
assign cj_6144[6107] = cin[2269];
assign cj_6144[6108] = cin[4356];
assign cj_6144[6109] = cin[1259];
assign cj_6144[6110] = cin[5266];
assign cj_6144[6111] = cin[4089];
assign cj_6144[6112] = cin[3872];
assign cj_6144[6113] = cin[4615];
assign cj_6144[6114] = cin[174];
assign cj_6144[6115] = cin[2837];
assign cj_6144[6116] = cin[316];
assign cj_6144[6117] = cin[4899];
assign cj_6144[6118] = cin[4298];
assign cj_6144[6119] = cin[4657];
assign cj_6144[6120] = cin[5976];
assign cj_6144[6121] = cin[2111];
assign cj_6144[6122] = cin[5350];
assign cj_6144[6123] = cin[3405];
assign cj_6144[6124] = cin[2420];
assign cj_6144[6125] = cin[2395];
assign cj_6144[6126] = cin[3330];
assign cj_6144[6127] = cin[5225];
assign cj_6144[6128] = cin[1936];
assign cj_6144[6129] = cin[5751];
assign cj_6144[6130] = cin[4382];
assign cj_6144[6131] = cin[3973];
assign cj_6144[6132] = cin[4524];
assign cj_6144[6133] = cin[6035];
assign cj_6144[6134] = cin[2362];
assign cj_6144[6135] = cin[5793];
assign cj_6144[6136] = cin[4040];
assign cj_6144[6137] = cin[3247];
assign cj_6144[6138] = cin[3414];
assign cj_6144[6139] = cin[4541];
assign cj_6144[6140] = cin[484];
assign cj_6144[6141] = cin[3531];
assign cj_6144[6142] = cin[1394];
assign cj_6144[6143] = cin[217];






endmodule

`endif