`ifndef CODER_INTERLEAVER_H
`define CODER_INTERLEAVER_H

module coder_interleaver (
	input [6143:0] cin,    // Clock
	input K_eq_6144,
	output [6143:0] cout,
	output [6143:0] ciout
);
	
	//c pi i wires given k
	wire [6143:0] cj_6144, cj_1056;

	//ci wires
	wire [6143:0] ci_6144;
	wire [1055:0] ci_1056;

	assign ci_6144 = cin;

	assign ciout = K_eq_6144?ci_6144:{5088'b0,ci_1056};

	//assigned in loops

	parameter f1_6144=263;

	parameter f1_1056=17;

	parameter f2_6144=480;

	parameter f2_1056=66;

	//for j from 0 to 6143
	genvar  j;
	generate
		for (j=0;j<4800;j=j+1)
		begin: loop0to4799
			assign cout[j]=K_eq_6144?cj_6144[j]:cj_1056[j];

		end
	endgenerate

	//for j2 from 0 to 6143
	genvar  j2;
	generate
		for (j2=4800;j2<6144;j2=j2+1)
		begin: loop4800to6143
			assign cout[j2]=K_eq_6144?cj_6144[j2]:cj_1056[j2];
		end
	endgenerate

	//for j from 0 to 1055

	// cj_6144[j]=cin[(f1_6144*j+f2_6144*j*j)%6144]

	// cj_1056[j]=cin[(f1_1056*j+f2_1056*j*j)%1056]

	genvar  i1;
	generate
		for (i1=0;i1<1056;i1=i1+1)
		begin: loop0to1055
			assign cj_6144[i1]=ci_6144[(f1_6144*i1+f2_6144*i1*i1) % 6144];
			assign cj_1056[i1]=ci_1056[(f1_1056*i1+f2_1056*i1*i1) % 1056];
			
			//no particular reason added here
			// to achieve: assign ci_6144 = cin[0:6143];
			//				&assign ci_1056 = cin[5088:6143];
			//assign ci_6144[i1] = cin[6143-i1];
			assign ci_1056[i1] = cin[5088+i1];
		end
	endgenerate


	//for j from 1056 to 2100
	genvar  i2;
	generate
		for (i2=1056;i2<2100;i2=i2+1)
		begin: loop1056to2099
			assign cj_6144[i2]=ci_6144[(f1_6144*i2+f2_6144*i2*i2)%6144];
			assign cj_1056[i2]=1'b0;

			//no particular reason added here
			// to achieve: assign ci_6144 = cin[0:6143];
			//assign ci_6144[i2] = cin[6143-i2];
		end
	endgenerate

	genvar  i3;
	generate
		for (i3=2100;i3<6144;i3=i3+1)
		begin: loop2100to6144
			//assign cj_6144[i3]=cin[(f1_6144*i3+f2_6144*i3*i3)%6144];
			assign cj_1056[i3]=1'b0;

			//no particular reason added here
			// to achieve: assign ci_6144 = cin[0:6143];
			//assign ci_6144[i3] = cin[6143-i3];
		end
	endgenerate


	assign cj_6144[2100] = ci_6144[876];
	assign cj_6144[2101] = ci_6144[2387];
	assign cj_6144[2102] = ci_6144[4858];
	assign cj_6144[2103] = ci_6144[2145];
	assign cj_6144[2104] = ci_6144[392];
	assign cj_6144[2105] = ci_6144[5743];
	assign cj_6144[2106] = ci_6144[5910];
	assign cj_6144[2107] = ci_6144[893];
	assign cj_6144[2108] = ci_6144[2980];
	assign cj_6144[2109] = ci_6144[6027];
	assign cj_6144[2110] = ci_6144[3890];
	assign cj_6144[2111] = ci_6144[2713];
	assign cj_6144[2112] = ci_6144[2496];
	assign cj_6144[2113] = ci_6144[3239];
	assign cj_6144[2114] = ci_6144[4942];
	assign cj_6144[2115] = ci_6144[1461];
	assign cj_6144[2116] = ci_6144[5084];
	assign cj_6144[2117] = ci_6144[3523];
	assign cj_6144[2118] = ci_6144[2922];
	assign cj_6144[2119] = ci_6144[3281];
	assign cj_6144[2120] = ci_6144[4600];
	assign cj_6144[2121] = ci_6144[735];
	assign cj_6144[2122] = ci_6144[3974];
	assign cj_6144[2123] = ci_6144[2029];
	assign cj_6144[2124] = ci_6144[1044];
	assign cj_6144[2125] = ci_6144[1019];
	assign cj_6144[2126] = ci_6144[1954];
	assign cj_6144[2127] = ci_6144[3849];
	assign cj_6144[2128] = ci_6144[560];
	assign cj_6144[2129] = ci_6144[4375];
	assign cj_6144[2130] = ci_6144[3006];
	assign cj_6144[2131] = ci_6144[2597];
	assign cj_6144[2132] = ci_6144[3148];
	assign cj_6144[2133] = ci_6144[4659];
	assign cj_6144[2134] = ci_6144[986];
	assign cj_6144[2135] = ci_6144[4417];
	assign cj_6144[2136] = ci_6144[2664];
	assign cj_6144[2137] = ci_6144[1871];
	assign cj_6144[2138] = ci_6144[2038];
	assign cj_6144[2139] = ci_6144[3165];
	assign cj_6144[2140] = ci_6144[5252];
	assign cj_6144[2141] = ci_6144[2155];
	assign cj_6144[2142] = ci_6144[18];
	assign cj_6144[2143] = ci_6144[4985];
	assign cj_6144[2144] = ci_6144[4768];
	assign cj_6144[2145] = ci_6144[5511];
	assign cj_6144[2146] = ci_6144[1070];
	assign cj_6144[2147] = ci_6144[3733];
	assign cj_6144[2148] = ci_6144[1212];
	assign cj_6144[2149] = ci_6144[5795];
	assign cj_6144[2150] = ci_6144[5194];
	assign cj_6144[2151] = ci_6144[5553];
	assign cj_6144[2152] = ci_6144[728];
	assign cj_6144[2153] = ci_6144[3007];
	assign cj_6144[2154] = ci_6144[102];
	assign cj_6144[2155] = ci_6144[4301];
	assign cj_6144[2156] = ci_6144[3316];
	assign cj_6144[2157] = ci_6144[3291];
	assign cj_6144[2158] = ci_6144[4226];
	assign cj_6144[2159] = ci_6144[6121];
	assign cj_6144[2160] = ci_6144[2832];
	assign cj_6144[2161] = ci_6144[503];
	assign cj_6144[2162] = ci_6144[5278];
	assign cj_6144[2163] = ci_6144[4869];
	assign cj_6144[2164] = ci_6144[5420];
	assign cj_6144[2165] = ci_6144[787];
	assign cj_6144[2166] = ci_6144[3258];
	assign cj_6144[2167] = ci_6144[545];
	assign cj_6144[2168] = ci_6144[4936];
	assign cj_6144[2169] = ci_6144[4143];
	assign cj_6144[2170] = ci_6144[4310];
	assign cj_6144[2171] = ci_6144[5437];
	assign cj_6144[2172] = ci_6144[1380];
	assign cj_6144[2173] = ci_6144[4427];
	assign cj_6144[2174] = ci_6144[2290];
	assign cj_6144[2175] = ci_6144[1113];
	assign cj_6144[2176] = ci_6144[896];
	assign cj_6144[2177] = ci_6144[1639];
	assign cj_6144[2178] = ci_6144[3342];
	assign cj_6144[2179] = ci_6144[6005];
	assign cj_6144[2180] = ci_6144[3484];
	assign cj_6144[2181] = ci_6144[1923];
	assign cj_6144[2182] = ci_6144[1322];
	assign cj_6144[2183] = ci_6144[1681];
	assign cj_6144[2184] = ci_6144[3000];
	assign cj_6144[2185] = ci_6144[5279];
	assign cj_6144[2186] = ci_6144[2374];
	assign cj_6144[2187] = ci_6144[429];
	assign cj_6144[2188] = ci_6144[5588];
	assign cj_6144[2189] = ci_6144[5563];
	assign cj_6144[2190] = ci_6144[354];
	assign cj_6144[2191] = ci_6144[2249];
	assign cj_6144[2192] = ci_6144[5104];
	assign cj_6144[2193] = ci_6144[2775];
	assign cj_6144[2194] = ci_6144[1406];
	assign cj_6144[2195] = ci_6144[997];
	assign cj_6144[2196] = ci_6144[1548];
	assign cj_6144[2197] = ci_6144[3059];
	assign cj_6144[2198] = ci_6144[5530];
	assign cj_6144[2199] = ci_6144[2817];
	assign cj_6144[2200] = ci_6144[1064];
	assign cj_6144[2201] = ci_6144[271];
	assign cj_6144[2202] = ci_6144[438];
	assign cj_6144[2203] = ci_6144[1565];
	assign cj_6144[2204] = ci_6144[3652];
	assign cj_6144[2205] = ci_6144[555];
	assign cj_6144[2206] = ci_6144[4562];
	assign cj_6144[2207] = ci_6144[3385];
	assign cj_6144[2208] = ci_6144[3168];
	assign cj_6144[2209] = ci_6144[3911];
	assign cj_6144[2210] = ci_6144[5614];
	assign cj_6144[2211] = ci_6144[2133];
	assign cj_6144[2212] = ci_6144[5756];
	assign cj_6144[2213] = ci_6144[4195];
	assign cj_6144[2214] = ci_6144[3594];
	assign cj_6144[2215] = ci_6144[3953];
	assign cj_6144[2216] = ci_6144[5272];
	assign cj_6144[2217] = ci_6144[1407];
	assign cj_6144[2218] = ci_6144[4646];
	assign cj_6144[2219] = ci_6144[2701];
	assign cj_6144[2220] = ci_6144[1716];
	assign cj_6144[2221] = ci_6144[1691];
	assign cj_6144[2222] = ci_6144[2626];
	assign cj_6144[2223] = ci_6144[4521];
	assign cj_6144[2224] = ci_6144[1232];
	assign cj_6144[2225] = ci_6144[5047];
	assign cj_6144[2226] = ci_6144[3678];
	assign cj_6144[2227] = ci_6144[3269];
	assign cj_6144[2228] = ci_6144[3820];
	assign cj_6144[2229] = ci_6144[5331];
	assign cj_6144[2230] = ci_6144[1658];
	assign cj_6144[2231] = ci_6144[5089];
	assign cj_6144[2232] = ci_6144[3336];
	assign cj_6144[2233] = ci_6144[2543];
	assign cj_6144[2234] = ci_6144[2710];
	assign cj_6144[2235] = ci_6144[3837];
	assign cj_6144[2236] = ci_6144[5924];
	assign cj_6144[2237] = ci_6144[2827];
	assign cj_6144[2238] = ci_6144[690];
	assign cj_6144[2239] = ci_6144[5657];
	assign cj_6144[2240] = ci_6144[5440];
	assign cj_6144[2241] = ci_6144[39];
	assign cj_6144[2242] = ci_6144[1742];
	assign cj_6144[2243] = ci_6144[4405];
	assign cj_6144[2244] = ci_6144[1884];
	assign cj_6144[2245] = ci_6144[323];
	assign cj_6144[2246] = ci_6144[5866];
	assign cj_6144[2247] = ci_6144[81];
	assign cj_6144[2248] = ci_6144[1400];
	assign cj_6144[2249] = ci_6144[3679];
	assign cj_6144[2250] = ci_6144[774];
	assign cj_6144[2251] = ci_6144[4973];
	assign cj_6144[2252] = ci_6144[3988];
	assign cj_6144[2253] = ci_6144[3963];
	assign cj_6144[2254] = ci_6144[4898];
	assign cj_6144[2255] = ci_6144[649];
	assign cj_6144[2256] = ci_6144[3504];
	assign cj_6144[2257] = ci_6144[1175];
	assign cj_6144[2258] = ci_6144[5950];
	assign cj_6144[2259] = ci_6144[5541];
	assign cj_6144[2260] = ci_6144[6092];
	assign cj_6144[2261] = ci_6144[1459];
	assign cj_6144[2262] = ci_6144[3930];
	assign cj_6144[2263] = ci_6144[1217];
	assign cj_6144[2264] = ci_6144[5608];
	assign cj_6144[2265] = ci_6144[4815];
	assign cj_6144[2266] = ci_6144[4982];
	assign cj_6144[2267] = ci_6144[6109];
	assign cj_6144[2268] = ci_6144[2052];
	assign cj_6144[2269] = ci_6144[5099];
	assign cj_6144[2270] = ci_6144[2962];
	assign cj_6144[2271] = ci_6144[1785];
	assign cj_6144[2272] = ci_6144[1568];
	assign cj_6144[2273] = ci_6144[2311];
	assign cj_6144[2274] = ci_6144[4014];
	assign cj_6144[2275] = ci_6144[533];
	assign cj_6144[2276] = ci_6144[4156];
	assign cj_6144[2277] = ci_6144[2595];
	assign cj_6144[2278] = ci_6144[1994];
	assign cj_6144[2279] = ci_6144[2353];
	assign cj_6144[2280] = ci_6144[3672];
	assign cj_6144[2281] = ci_6144[5951];
	assign cj_6144[2282] = ci_6144[3046];
	assign cj_6144[2283] = ci_6144[1101];
	assign cj_6144[2284] = ci_6144[116];
	assign cj_6144[2285] = ci_6144[91];
	assign cj_6144[2286] = ci_6144[1026];
	assign cj_6144[2287] = ci_6144[2921];
	assign cj_6144[2288] = ci_6144[5776];
	assign cj_6144[2289] = ci_6144[3447];
	assign cj_6144[2290] = ci_6144[2078];
	assign cj_6144[2291] = ci_6144[1669];
	assign cj_6144[2292] = ci_6144[2220];
	assign cj_6144[2293] = ci_6144[3731];
	assign cj_6144[2294] = ci_6144[58];
	assign cj_6144[2295] = ci_6144[3489];
	assign cj_6144[2296] = ci_6144[1736];
	assign cj_6144[2297] = ci_6144[943];
	assign cj_6144[2298] = ci_6144[1110];
	assign cj_6144[2299] = ci_6144[2237];
	assign cj_6144[2300] = ci_6144[4324];
	assign cj_6144[2301] = ci_6144[1227];
	assign cj_6144[2302] = ci_6144[5234];
	assign cj_6144[2303] = ci_6144[4057];
	assign cj_6144[2304] = ci_6144[3840];
	assign cj_6144[2305] = ci_6144[4583];
	assign cj_6144[2306] = ci_6144[142];
	assign cj_6144[2307] = ci_6144[2805];
	assign cj_6144[2308] = ci_6144[284];
	assign cj_6144[2309] = ci_6144[4867];
	assign cj_6144[2310] = ci_6144[4266];
	assign cj_6144[2311] = ci_6144[4625];
	assign cj_6144[2312] = ci_6144[5944];
	assign cj_6144[2313] = ci_6144[2079];
	assign cj_6144[2314] = ci_6144[5318];
	assign cj_6144[2315] = ci_6144[3373];
	assign cj_6144[2316] = ci_6144[2388];
	assign cj_6144[2317] = ci_6144[2363];
	assign cj_6144[2318] = ci_6144[3298];
	assign cj_6144[2319] = ci_6144[5193];
	assign cj_6144[2320] = ci_6144[1904];
	assign cj_6144[2321] = ci_6144[5719];
	assign cj_6144[2322] = ci_6144[4350];
	assign cj_6144[2323] = ci_6144[3941];
	assign cj_6144[2324] = ci_6144[4492];
	assign cj_6144[2325] = ci_6144[6003];
	assign cj_6144[2326] = ci_6144[2330];
	assign cj_6144[2327] = ci_6144[5761];
	assign cj_6144[2328] = ci_6144[4008];
	assign cj_6144[2329] = ci_6144[3215];
	assign cj_6144[2330] = ci_6144[3382];
	assign cj_6144[2331] = ci_6144[4509];
	assign cj_6144[2332] = ci_6144[452];
	assign cj_6144[2333] = ci_6144[3499];
	assign cj_6144[2334] = ci_6144[1362];
	assign cj_6144[2335] = ci_6144[185];
	assign cj_6144[2336] = ci_6144[6112];
	assign cj_6144[2337] = ci_6144[711];
	assign cj_6144[2338] = ci_6144[2414];
	assign cj_6144[2339] = ci_6144[5077];
	assign cj_6144[2340] = ci_6144[2556];
	assign cj_6144[2341] = ci_6144[995];
	assign cj_6144[2342] = ci_6144[394];
	assign cj_6144[2343] = ci_6144[753];
	assign cj_6144[2344] = ci_6144[2072];
	assign cj_6144[2345] = ci_6144[4351];
	assign cj_6144[2346] = ci_6144[1446];
	assign cj_6144[2347] = ci_6144[5645];
	assign cj_6144[2348] = ci_6144[4660];
	assign cj_6144[2349] = ci_6144[4635];
	assign cj_6144[2350] = ci_6144[5570];
	assign cj_6144[2351] = ci_6144[1321];
	assign cj_6144[2352] = ci_6144[4176];
	assign cj_6144[2353] = ci_6144[1847];
	assign cj_6144[2354] = ci_6144[478];
	assign cj_6144[2355] = ci_6144[69];
	assign cj_6144[2356] = ci_6144[620];
	assign cj_6144[2357] = ci_6144[2131];
	assign cj_6144[2358] = ci_6144[4602];
	assign cj_6144[2359] = ci_6144[1889];
	assign cj_6144[2360] = ci_6144[136];
	assign cj_6144[2361] = ci_6144[5487];
	assign cj_6144[2362] = ci_6144[5654];
	assign cj_6144[2363] = ci_6144[637];
	assign cj_6144[2364] = ci_6144[2724];
	assign cj_6144[2365] = ci_6144[5771];
	assign cj_6144[2366] = ci_6144[3634];
	assign cj_6144[2367] = ci_6144[2457];
	assign cj_6144[2368] = ci_6144[2240];
	assign cj_6144[2369] = ci_6144[2983];
	assign cj_6144[2370] = ci_6144[4686];
	assign cj_6144[2371] = ci_6144[1205];
	assign cj_6144[2372] = ci_6144[4828];
	assign cj_6144[2373] = ci_6144[3267];
	assign cj_6144[2374] = ci_6144[2666];
	assign cj_6144[2375] = ci_6144[3025];
	assign cj_6144[2376] = ci_6144[4344];
	assign cj_6144[2377] = ci_6144[479];
	assign cj_6144[2378] = ci_6144[3718];
	assign cj_6144[2379] = ci_6144[1773];
	assign cj_6144[2380] = ci_6144[788];
	assign cj_6144[2381] = ci_6144[763];
	assign cj_6144[2382] = ci_6144[1698];
	assign cj_6144[2383] = ci_6144[3593];
	assign cj_6144[2384] = ci_6144[304];
	assign cj_6144[2385] = ci_6144[4119];
	assign cj_6144[2386] = ci_6144[2750];
	assign cj_6144[2387] = ci_6144[2341];
	assign cj_6144[2388] = ci_6144[2892];
	assign cj_6144[2389] = ci_6144[4403];
	assign cj_6144[2390] = ci_6144[730];
	assign cj_6144[2391] = ci_6144[4161];
	assign cj_6144[2392] = ci_6144[2408];
	assign cj_6144[2393] = ci_6144[1615];
	assign cj_6144[2394] = ci_6144[1782];
	assign cj_6144[2395] = ci_6144[2909];
	assign cj_6144[2396] = ci_6144[4996];
	assign cj_6144[2397] = ci_6144[1899];
	assign cj_6144[2398] = ci_6144[5906];
	assign cj_6144[2399] = ci_6144[4729];
	assign cj_6144[2400] = ci_6144[4512];
	assign cj_6144[2401] = ci_6144[5255];
	assign cj_6144[2402] = ci_6144[814];
	assign cj_6144[2403] = ci_6144[3477];
	assign cj_6144[2404] = ci_6144[956];
	assign cj_6144[2405] = ci_6144[5539];
	assign cj_6144[2406] = ci_6144[4938];
	assign cj_6144[2407] = ci_6144[5297];
	assign cj_6144[2408] = ci_6144[472];
	assign cj_6144[2409] = ci_6144[2751];
	assign cj_6144[2410] = ci_6144[5990];
	assign cj_6144[2411] = ci_6144[4045];
	assign cj_6144[2412] = ci_6144[3060];
	assign cj_6144[2413] = ci_6144[3035];
	assign cj_6144[2414] = ci_6144[3970];
	assign cj_6144[2415] = ci_6144[5865];
	assign cj_6144[2416] = ci_6144[2576];
	assign cj_6144[2417] = ci_6144[247];
	assign cj_6144[2418] = ci_6144[5022];
	assign cj_6144[2419] = ci_6144[4613];
	assign cj_6144[2420] = ci_6144[5164];
	assign cj_6144[2421] = ci_6144[531];
	assign cj_6144[2422] = ci_6144[3002];
	assign cj_6144[2423] = ci_6144[289];
	assign cj_6144[2424] = ci_6144[4680];
	assign cj_6144[2425] = ci_6144[3887];
	assign cj_6144[2426] = ci_6144[4054];
	assign cj_6144[2427] = ci_6144[5181];
	assign cj_6144[2428] = ci_6144[1124];
	assign cj_6144[2429] = ci_6144[4171];
	assign cj_6144[2430] = ci_6144[2034];
	assign cj_6144[2431] = ci_6144[857];
	assign cj_6144[2432] = ci_6144[640];
	assign cj_6144[2433] = ci_6144[1383];
	assign cj_6144[2434] = ci_6144[3086];
	assign cj_6144[2435] = ci_6144[5749];
	assign cj_6144[2436] = ci_6144[3228];
	assign cj_6144[2437] = ci_6144[1667];
	assign cj_6144[2438] = ci_6144[1066];
	assign cj_6144[2439] = ci_6144[1425];
	assign cj_6144[2440] = ci_6144[2744];
	assign cj_6144[2441] = ci_6144[5023];
	assign cj_6144[2442] = ci_6144[2118];
	assign cj_6144[2443] = ci_6144[173];
	assign cj_6144[2444] = ci_6144[5332];
	assign cj_6144[2445] = ci_6144[5307];
	assign cj_6144[2446] = ci_6144[98];
	assign cj_6144[2447] = ci_6144[1993];
	assign cj_6144[2448] = ci_6144[4848];
	assign cj_6144[2449] = ci_6144[2519];
	assign cj_6144[2450] = ci_6144[1150];
	assign cj_6144[2451] = ci_6144[741];
	assign cj_6144[2452] = ci_6144[1292];
	assign cj_6144[2453] = ci_6144[2803];
	assign cj_6144[2454] = ci_6144[5274];
	assign cj_6144[2455] = ci_6144[2561];
	assign cj_6144[2456] = ci_6144[808];
	assign cj_6144[2457] = ci_6144[15];
	assign cj_6144[2458] = ci_6144[182];
	assign cj_6144[2459] = ci_6144[1309];
	assign cj_6144[2460] = ci_6144[3396];
	assign cj_6144[2461] = ci_6144[299];
	assign cj_6144[2462] = ci_6144[4306];
	assign cj_6144[2463] = ci_6144[3129];
	assign cj_6144[2464] = ci_6144[2912];
	assign cj_6144[2465] = ci_6144[3655];
	assign cj_6144[2466] = ci_6144[5358];
	assign cj_6144[2467] = ci_6144[1877];
	assign cj_6144[2468] = ci_6144[5500];
	assign cj_6144[2469] = ci_6144[3939];
	assign cj_6144[2470] = ci_6144[3338];
	assign cj_6144[2471] = ci_6144[3697];
	assign cj_6144[2472] = ci_6144[5016];
	assign cj_6144[2473] = ci_6144[1151];
	assign cj_6144[2474] = ci_6144[4390];
	assign cj_6144[2475] = ci_6144[2445];
	assign cj_6144[2476] = ci_6144[1460];
	assign cj_6144[2477] = ci_6144[1435];
	assign cj_6144[2478] = ci_6144[2370];
	assign cj_6144[2479] = ci_6144[4265];
	assign cj_6144[2480] = ci_6144[976];
	assign cj_6144[2481] = ci_6144[4791];
	assign cj_6144[2482] = ci_6144[3422];
	assign cj_6144[2483] = ci_6144[3013];
	assign cj_6144[2484] = ci_6144[3564];
	assign cj_6144[2485] = ci_6144[5075];
	assign cj_6144[2486] = ci_6144[1402];
	assign cj_6144[2487] = ci_6144[4833];
	assign cj_6144[2488] = ci_6144[3080];
	assign cj_6144[2489] = ci_6144[2287];
	assign cj_6144[2490] = ci_6144[2454];
	assign cj_6144[2491] = ci_6144[3581];
	assign cj_6144[2492] = ci_6144[5668];
	assign cj_6144[2493] = ci_6144[2571];
	assign cj_6144[2494] = ci_6144[434];
	assign cj_6144[2495] = ci_6144[5401];
	assign cj_6144[2496] = ci_6144[5184];
	assign cj_6144[2497] = ci_6144[5927];
	assign cj_6144[2498] = ci_6144[1486];
	assign cj_6144[2499] = ci_6144[4149];
	assign cj_6144[2500] = ci_6144[1628];
	assign cj_6144[2501] = ci_6144[67];
	assign cj_6144[2502] = ci_6144[5610];
	assign cj_6144[2503] = ci_6144[5969];
	assign cj_6144[2504] = ci_6144[1144];
	assign cj_6144[2505] = ci_6144[3423];
	assign cj_6144[2506] = ci_6144[518];
	assign cj_6144[2507] = ci_6144[4717];
	assign cj_6144[2508] = ci_6144[3732];
	assign cj_6144[2509] = ci_6144[3707];
	assign cj_6144[2510] = ci_6144[4642];
	assign cj_6144[2511] = ci_6144[393];
	assign cj_6144[2512] = ci_6144[3248];
	assign cj_6144[2513] = ci_6144[919];
	assign cj_6144[2514] = ci_6144[5694];
	assign cj_6144[2515] = ci_6144[5285];
	assign cj_6144[2516] = ci_6144[5836];
	assign cj_6144[2517] = ci_6144[1203];
	assign cj_6144[2518] = ci_6144[3674];
	assign cj_6144[2519] = ci_6144[961];
	assign cj_6144[2520] = ci_6144[5352];
	assign cj_6144[2521] = ci_6144[4559];
	assign cj_6144[2522] = ci_6144[4726];
	assign cj_6144[2523] = ci_6144[5853];
	assign cj_6144[2524] = ci_6144[1796];
	assign cj_6144[2525] = ci_6144[4843];
	assign cj_6144[2526] = ci_6144[2706];
	assign cj_6144[2527] = ci_6144[1529];
	assign cj_6144[2528] = ci_6144[1312];
	assign cj_6144[2529] = ci_6144[2055];
	assign cj_6144[2530] = ci_6144[3758];
	assign cj_6144[2531] = ci_6144[277];
	assign cj_6144[2532] = ci_6144[3900];
	assign cj_6144[2533] = ci_6144[2339];
	assign cj_6144[2534] = ci_6144[1738];
	assign cj_6144[2535] = ci_6144[2097];
	assign cj_6144[2536] = ci_6144[3416];
	assign cj_6144[2537] = ci_6144[5695];
	assign cj_6144[2538] = ci_6144[2790];
	assign cj_6144[2539] = ci_6144[845];
	assign cj_6144[2540] = ci_6144[6004];
	assign cj_6144[2541] = ci_6144[5979];
	assign cj_6144[2542] = ci_6144[770];
	assign cj_6144[2543] = ci_6144[2665];
	assign cj_6144[2544] = ci_6144[5520];
	assign cj_6144[2545] = ci_6144[3191];
	assign cj_6144[2546] = ci_6144[1822];
	assign cj_6144[2547] = ci_6144[1413];
	assign cj_6144[2548] = ci_6144[1964];
	assign cj_6144[2549] = ci_6144[3475];
	assign cj_6144[2550] = ci_6144[5946];
	assign cj_6144[2551] = ci_6144[3233];
	assign cj_6144[2552] = ci_6144[1480];
	assign cj_6144[2553] = ci_6144[687];
	assign cj_6144[2554] = ci_6144[854];
	assign cj_6144[2555] = ci_6144[1981];
	assign cj_6144[2556] = ci_6144[4068];
	assign cj_6144[2557] = ci_6144[971];
	assign cj_6144[2558] = ci_6144[4978];
	assign cj_6144[2559] = ci_6144[3801];
	assign cj_6144[2560] = ci_6144[3584];
	assign cj_6144[2561] = ci_6144[4327];
	assign cj_6144[2562] = ci_6144[6030];
	assign cj_6144[2563] = ci_6144[2549];
	assign cj_6144[2564] = ci_6144[28];
	assign cj_6144[2565] = ci_6144[4611];
	assign cj_6144[2566] = ci_6144[4010];
	assign cj_6144[2567] = ci_6144[4369];
	assign cj_6144[2568] = ci_6144[5688];
	assign cj_6144[2569] = ci_6144[1823];
	assign cj_6144[2570] = ci_6144[5062];
	assign cj_6144[2571] = ci_6144[3117];
	assign cj_6144[2572] = ci_6144[2132];
	assign cj_6144[2573] = ci_6144[2107];
	assign cj_6144[2574] = ci_6144[3042];
	assign cj_6144[2575] = ci_6144[4937];
	assign cj_6144[2576] = ci_6144[1648];
	assign cj_6144[2577] = ci_6144[5463];
	assign cj_6144[2578] = ci_6144[4094];
	assign cj_6144[2579] = ci_6144[3685];
	assign cj_6144[2580] = ci_6144[4236];
	assign cj_6144[2581] = ci_6144[5747];
	assign cj_6144[2582] = ci_6144[2074];
	assign cj_6144[2583] = ci_6144[5505];
	assign cj_6144[2584] = ci_6144[3752];
	assign cj_6144[2585] = ci_6144[2959];
	assign cj_6144[2586] = ci_6144[3126];
	assign cj_6144[2587] = ci_6144[4253];
	assign cj_6144[2588] = ci_6144[196];
	assign cj_6144[2589] = ci_6144[3243];
	assign cj_6144[2590] = ci_6144[1106];
	assign cj_6144[2591] = ci_6144[6073];
	assign cj_6144[2592] = ci_6144[5856];
	assign cj_6144[2593] = ci_6144[455];
	assign cj_6144[2594] = ci_6144[2158];
	assign cj_6144[2595] = ci_6144[4821];
	assign cj_6144[2596] = ci_6144[2300];
	assign cj_6144[2597] = ci_6144[739];
	assign cj_6144[2598] = ci_6144[138];
	assign cj_6144[2599] = ci_6144[497];
	assign cj_6144[2600] = ci_6144[1816];
	assign cj_6144[2601] = ci_6144[4095];
	assign cj_6144[2602] = ci_6144[1190];
	assign cj_6144[2603] = ci_6144[5389];
	assign cj_6144[2604] = ci_6144[4404];
	assign cj_6144[2605] = ci_6144[4379];
	assign cj_6144[2606] = ci_6144[5314];
	assign cj_6144[2607] = ci_6144[1065];
	assign cj_6144[2608] = ci_6144[3920];
	assign cj_6144[2609] = ci_6144[1591];
	assign cj_6144[2610] = ci_6144[222];
	assign cj_6144[2611] = ci_6144[5957];
	assign cj_6144[2612] = ci_6144[364];
	assign cj_6144[2613] = ci_6144[1875];
	assign cj_6144[2614] = ci_6144[4346];
	assign cj_6144[2615] = ci_6144[1633];
	assign cj_6144[2616] = ci_6144[6024];
	assign cj_6144[2617] = ci_6144[5231];
	assign cj_6144[2618] = ci_6144[5398];
	assign cj_6144[2619] = ci_6144[381];
	assign cj_6144[2620] = ci_6144[2468];
	assign cj_6144[2621] = ci_6144[5515];
	assign cj_6144[2622] = ci_6144[3378];
	assign cj_6144[2623] = ci_6144[2201];
	assign cj_6144[2624] = ci_6144[1984];
	assign cj_6144[2625] = ci_6144[2727];
	assign cj_6144[2626] = ci_6144[4430];
	assign cj_6144[2627] = ci_6144[949];
	assign cj_6144[2628] = ci_6144[4572];
	assign cj_6144[2629] = ci_6144[3011];
	assign cj_6144[2630] = ci_6144[2410];
	assign cj_6144[2631] = ci_6144[2769];
	assign cj_6144[2632] = ci_6144[4088];
	assign cj_6144[2633] = ci_6144[223];
	assign cj_6144[2634] = ci_6144[3462];
	assign cj_6144[2635] = ci_6144[1517];
	assign cj_6144[2636] = ci_6144[532];
	assign cj_6144[2637] = ci_6144[507];
	assign cj_6144[2638] = ci_6144[1442];
	assign cj_6144[2639] = ci_6144[3337];
	assign cj_6144[2640] = ci_6144[48];
	assign cj_6144[2641] = ci_6144[3863];
	assign cj_6144[2642] = ci_6144[2494];
	assign cj_6144[2643] = ci_6144[2085];
	assign cj_6144[2644] = ci_6144[2636];
	assign cj_6144[2645] = ci_6144[4147];
	assign cj_6144[2646] = ci_6144[474];
	assign cj_6144[2647] = ci_6144[3905];
	assign cj_6144[2648] = ci_6144[2152];
	assign cj_6144[2649] = ci_6144[1359];
	assign cj_6144[2650] = ci_6144[1526];
	assign cj_6144[2651] = ci_6144[2653];
	assign cj_6144[2652] = ci_6144[4740];
	assign cj_6144[2653] = ci_6144[1643];
	assign cj_6144[2654] = ci_6144[5650];
	assign cj_6144[2655] = ci_6144[4473];
	assign cj_6144[2656] = ci_6144[4256];
	assign cj_6144[2657] = ci_6144[4999];
	assign cj_6144[2658] = ci_6144[558];
	assign cj_6144[2659] = ci_6144[3221];
	assign cj_6144[2660] = ci_6144[700];
	assign cj_6144[2661] = ci_6144[5283];
	assign cj_6144[2662] = ci_6144[4682];
	assign cj_6144[2663] = ci_6144[5041];
	assign cj_6144[2664] = ci_6144[216];
	assign cj_6144[2665] = ci_6144[2495];
	assign cj_6144[2666] = ci_6144[5734];
	assign cj_6144[2667] = ci_6144[3789];
	assign cj_6144[2668] = ci_6144[2804];
	assign cj_6144[2669] = ci_6144[2779];
	assign cj_6144[2670] = ci_6144[3714];
	assign cj_6144[2671] = ci_6144[5609];
	assign cj_6144[2672] = ci_6144[2320];
	assign cj_6144[2673] = ci_6144[6135];
	assign cj_6144[2674] = ci_6144[4766];
	assign cj_6144[2675] = ci_6144[4357];
	assign cj_6144[2676] = ci_6144[4908];
	assign cj_6144[2677] = ci_6144[275];
	assign cj_6144[2678] = ci_6144[2746];
	assign cj_6144[2679] = ci_6144[33];
	assign cj_6144[2680] = ci_6144[4424];
	assign cj_6144[2681] = ci_6144[3631];
	assign cj_6144[2682] = ci_6144[3798];
	assign cj_6144[2683] = ci_6144[4925];
	assign cj_6144[2684] = ci_6144[868];
	assign cj_6144[2685] = ci_6144[3915];
	assign cj_6144[2686] = ci_6144[1778];
	assign cj_6144[2687] = ci_6144[601];
	assign cj_6144[2688] = ci_6144[384];
	assign cj_6144[2689] = ci_6144[1127];
	assign cj_6144[2690] = ci_6144[2830];
	assign cj_6144[2691] = ci_6144[5493];
	assign cj_6144[2692] = ci_6144[2972];
	assign cj_6144[2693] = ci_6144[1411];
	assign cj_6144[2694] = ci_6144[810];
	assign cj_6144[2695] = ci_6144[1169];
	assign cj_6144[2696] = ci_6144[2488];
	assign cj_6144[2697] = ci_6144[4767];
	assign cj_6144[2698] = ci_6144[1862];
	assign cj_6144[2699] = ci_6144[6061];
	assign cj_6144[2700] = ci_6144[5076];
	assign cj_6144[2701] = ci_6144[5051];
	assign cj_6144[2702] = ci_6144[5986];
	assign cj_6144[2703] = ci_6144[1737];
	assign cj_6144[2704] = ci_6144[4592];
	assign cj_6144[2705] = ci_6144[2263];
	assign cj_6144[2706] = ci_6144[894];
	assign cj_6144[2707] = ci_6144[485];
	assign cj_6144[2708] = ci_6144[1036];
	assign cj_6144[2709] = ci_6144[2547];
	assign cj_6144[2710] = ci_6144[5018];
	assign cj_6144[2711] = ci_6144[2305];
	assign cj_6144[2712] = ci_6144[552];
	assign cj_6144[2713] = ci_6144[5903];
	assign cj_6144[2714] = ci_6144[6070];
	assign cj_6144[2715] = ci_6144[1053];
	assign cj_6144[2716] = ci_6144[3140];
	assign cj_6144[2717] = ci_6144[43];
	assign cj_6144[2718] = ci_6144[4050];
	assign cj_6144[2719] = ci_6144[2873];
	assign cj_6144[2720] = ci_6144[2656];
	assign cj_6144[2721] = ci_6144[3399];
	assign cj_6144[2722] = ci_6144[5102];
	assign cj_6144[2723] = ci_6144[1621];
	assign cj_6144[2724] = ci_6144[5244];
	assign cj_6144[2725] = ci_6144[3683];
	assign cj_6144[2726] = ci_6144[3082];
	assign cj_6144[2727] = ci_6144[3441];
	assign cj_6144[2728] = ci_6144[4760];
	assign cj_6144[2729] = ci_6144[895];
	assign cj_6144[2730] = ci_6144[4134];
	assign cj_6144[2731] = ci_6144[2189];
	assign cj_6144[2732] = ci_6144[1204];
	assign cj_6144[2733] = ci_6144[1179];
	assign cj_6144[2734] = ci_6144[2114];
	assign cj_6144[2735] = ci_6144[4009];
	assign cj_6144[2736] = ci_6144[720];
	assign cj_6144[2737] = ci_6144[4535];
	assign cj_6144[2738] = ci_6144[3166];
	assign cj_6144[2739] = ci_6144[2757];
	assign cj_6144[2740] = ci_6144[3308];
	assign cj_6144[2741] = ci_6144[4819];
	assign cj_6144[2742] = ci_6144[1146];
	assign cj_6144[2743] = ci_6144[4577];
	assign cj_6144[2744] = ci_6144[2824];
	assign cj_6144[2745] = ci_6144[2031];
	assign cj_6144[2746] = ci_6144[2198];
	assign cj_6144[2747] = ci_6144[3325];
	assign cj_6144[2748] = ci_6144[5412];
	assign cj_6144[2749] = ci_6144[2315];
	assign cj_6144[2750] = ci_6144[178];
	assign cj_6144[2751] = ci_6144[5145];
	assign cj_6144[2752] = ci_6144[4928];
	assign cj_6144[2753] = ci_6144[5671];
	assign cj_6144[2754] = ci_6144[1230];
	assign cj_6144[2755] = ci_6144[3893];
	assign cj_6144[2756] = ci_6144[1372];
	assign cj_6144[2757] = ci_6144[5955];
	assign cj_6144[2758] = ci_6144[5354];
	assign cj_6144[2759] = ci_6144[5713];
	assign cj_6144[2760] = ci_6144[888];
	assign cj_6144[2761] = ci_6144[3167];
	assign cj_6144[2762] = ci_6144[262];
	assign cj_6144[2763] = ci_6144[4461];
	assign cj_6144[2764] = ci_6144[3476];
	assign cj_6144[2765] = ci_6144[3451];
	assign cj_6144[2766] = ci_6144[4386];
	assign cj_6144[2767] = ci_6144[137];
	assign cj_6144[2768] = ci_6144[2992];
	assign cj_6144[2769] = ci_6144[663];
	assign cj_6144[2770] = ci_6144[5438];
	assign cj_6144[2771] = ci_6144[5029];
	assign cj_6144[2772] = ci_6144[5580];
	assign cj_6144[2773] = ci_6144[947];
	assign cj_6144[2774] = ci_6144[3418];
	assign cj_6144[2775] = ci_6144[705];
	assign cj_6144[2776] = ci_6144[5096];
	assign cj_6144[2777] = ci_6144[4303];
	assign cj_6144[2778] = ci_6144[4470];
	assign cj_6144[2779] = ci_6144[5597];
	assign cj_6144[2780] = ci_6144[1540];
	assign cj_6144[2781] = ci_6144[4587];
	assign cj_6144[2782] = ci_6144[2450];
	assign cj_6144[2783] = ci_6144[1273];
	assign cj_6144[2784] = ci_6144[1056];
	assign cj_6144[2785] = ci_6144[1799];
	assign cj_6144[2786] = ci_6144[3502];
	assign cj_6144[2787] = ci_6144[21];
	assign cj_6144[2788] = ci_6144[3644];
	assign cj_6144[2789] = ci_6144[2083];
	assign cj_6144[2790] = ci_6144[1482];
	assign cj_6144[2791] = ci_6144[1841];
	assign cj_6144[2792] = ci_6144[3160];
	assign cj_6144[2793] = ci_6144[5439];
	assign cj_6144[2794] = ci_6144[2534];
	assign cj_6144[2795] = ci_6144[589];
	assign cj_6144[2796] = ci_6144[5748];
	assign cj_6144[2797] = ci_6144[5723];
	assign cj_6144[2798] = ci_6144[514];
	assign cj_6144[2799] = ci_6144[2409];
	assign cj_6144[2800] = ci_6144[5264];
	assign cj_6144[2801] = ci_6144[2935];
	assign cj_6144[2802] = ci_6144[1566];
	assign cj_6144[2803] = ci_6144[1157];
	assign cj_6144[2804] = ci_6144[1708];
	assign cj_6144[2805] = ci_6144[3219];
	assign cj_6144[2806] = ci_6144[5690];
	assign cj_6144[2807] = ci_6144[2977];
	assign cj_6144[2808] = ci_6144[1224];
	assign cj_6144[2809] = ci_6144[431];
	assign cj_6144[2810] = ci_6144[598];
	assign cj_6144[2811] = ci_6144[1725];
	assign cj_6144[2812] = ci_6144[3812];
	assign cj_6144[2813] = ci_6144[715];
	assign cj_6144[2814] = ci_6144[4722];
	assign cj_6144[2815] = ci_6144[3545];
	assign cj_6144[2816] = ci_6144[3328];
	assign cj_6144[2817] = ci_6144[4071];
	assign cj_6144[2818] = ci_6144[5774];
	assign cj_6144[2819] = ci_6144[2293];
	assign cj_6144[2820] = ci_6144[5916];
	assign cj_6144[2821] = ci_6144[4355];
	assign cj_6144[2822] = ci_6144[3754];
	assign cj_6144[2823] = ci_6144[4113];
	assign cj_6144[2824] = ci_6144[5432];
	assign cj_6144[2825] = ci_6144[1567];
	assign cj_6144[2826] = ci_6144[4806];
	assign cj_6144[2827] = ci_6144[2861];
	assign cj_6144[2828] = ci_6144[1876];
	assign cj_6144[2829] = ci_6144[1851];
	assign cj_6144[2830] = ci_6144[2786];
	assign cj_6144[2831] = ci_6144[4681];
	assign cj_6144[2832] = ci_6144[1392];
	assign cj_6144[2833] = ci_6144[5207];
	assign cj_6144[2834] = ci_6144[3838];
	assign cj_6144[2835] = ci_6144[3429];
	assign cj_6144[2836] = ci_6144[3980];
	assign cj_6144[2837] = ci_6144[5491];
	assign cj_6144[2838] = ci_6144[1818];
	assign cj_6144[2839] = ci_6144[5249];
	assign cj_6144[2840] = ci_6144[3496];
	assign cj_6144[2841] = ci_6144[2703];
	assign cj_6144[2842] = ci_6144[2870];
	assign cj_6144[2843] = ci_6144[3997];
	assign cj_6144[2844] = ci_6144[6084];
	assign cj_6144[2845] = ci_6144[2987];
	assign cj_6144[2846] = ci_6144[850];
	assign cj_6144[2847] = ci_6144[5817];
	assign cj_6144[2848] = ci_6144[5600];
	assign cj_6144[2849] = ci_6144[199];
	assign cj_6144[2850] = ci_6144[1902];
	assign cj_6144[2851] = ci_6144[4565];
	assign cj_6144[2852] = ci_6144[2044];
	assign cj_6144[2853] = ci_6144[483];
	assign cj_6144[2854] = ci_6144[6026];
	assign cj_6144[2855] = ci_6144[241];
	assign cj_6144[2856] = ci_6144[1560];
	assign cj_6144[2857] = ci_6144[3839];
	assign cj_6144[2858] = ci_6144[934];
	assign cj_6144[2859] = ci_6144[5133];
	assign cj_6144[2860] = ci_6144[4148];
	assign cj_6144[2861] = ci_6144[4123];
	assign cj_6144[2862] = ci_6144[5058];
	assign cj_6144[2863] = ci_6144[809];
	assign cj_6144[2864] = ci_6144[3664];
	assign cj_6144[2865] = ci_6144[1335];
	assign cj_6144[2866] = ci_6144[6110];
	assign cj_6144[2867] = ci_6144[5701];
	assign cj_6144[2868] = ci_6144[108];
	assign cj_6144[2869] = ci_6144[1619];
	assign cj_6144[2870] = ci_6144[4090];
	assign cj_6144[2871] = ci_6144[1377];
	assign cj_6144[2872] = ci_6144[5768];
	assign cj_6144[2873] = ci_6144[4975];
	assign cj_6144[2874] = ci_6144[5142];
	assign cj_6144[2875] = ci_6144[125];
	assign cj_6144[2876] = ci_6144[2212];
	assign cj_6144[2877] = ci_6144[5259];
	assign cj_6144[2878] = ci_6144[3122];
	assign cj_6144[2879] = ci_6144[1945];
	assign cj_6144[2880] = ci_6144[1728];
	assign cj_6144[2881] = ci_6144[2471];
	assign cj_6144[2882] = ci_6144[4174];
	assign cj_6144[2883] = ci_6144[693];
	assign cj_6144[2884] = ci_6144[4316];
	assign cj_6144[2885] = ci_6144[2755];
	assign cj_6144[2886] = ci_6144[2154];
	assign cj_6144[2887] = ci_6144[2513];
	assign cj_6144[2888] = ci_6144[3832];
	assign cj_6144[2889] = ci_6144[6111];
	assign cj_6144[2890] = ci_6144[3206];
	assign cj_6144[2891] = ci_6144[1261];
	assign cj_6144[2892] = ci_6144[276];
	assign cj_6144[2893] = ci_6144[251];
	assign cj_6144[2894] = ci_6144[1186];
	assign cj_6144[2895] = ci_6144[3081];
	assign cj_6144[2896] = ci_6144[5936];
	assign cj_6144[2897] = ci_6144[3607];
	assign cj_6144[2898] = ci_6144[2238];
	assign cj_6144[2899] = ci_6144[1829];
	assign cj_6144[2900] = ci_6144[2380];
	assign cj_6144[2901] = ci_6144[3891];
	assign cj_6144[2902] = ci_6144[218];
	assign cj_6144[2903] = ci_6144[3649];
	assign cj_6144[2904] = ci_6144[1896];
	assign cj_6144[2905] = ci_6144[1103];
	assign cj_6144[2906] = ci_6144[1270];
	assign cj_6144[2907] = ci_6144[2397];
	assign cj_6144[2908] = ci_6144[4484];
	assign cj_6144[2909] = ci_6144[1387];
	assign cj_6144[2910] = ci_6144[5394];
	assign cj_6144[2911] = ci_6144[4217];
	assign cj_6144[2912] = ci_6144[4000];
	assign cj_6144[2913] = ci_6144[4743];
	assign cj_6144[2914] = ci_6144[302];
	assign cj_6144[2915] = ci_6144[2965];
	assign cj_6144[2916] = ci_6144[444];
	assign cj_6144[2917] = ci_6144[5027];
	assign cj_6144[2918] = ci_6144[4426];
	assign cj_6144[2919] = ci_6144[4785];
	assign cj_6144[2920] = ci_6144[6104];
	assign cj_6144[2921] = ci_6144[2239];
	assign cj_6144[2922] = ci_6144[5478];
	assign cj_6144[2923] = ci_6144[3533];
	assign cj_6144[2924] = ci_6144[2548];
	assign cj_6144[2925] = ci_6144[2523];
	assign cj_6144[2926] = ci_6144[3458];
	assign cj_6144[2927] = ci_6144[5353];
	assign cj_6144[2928] = ci_6144[2064];
	assign cj_6144[2929] = ci_6144[5879];
	assign cj_6144[2930] = ci_6144[4510];
	assign cj_6144[2931] = ci_6144[4101];
	assign cj_6144[2932] = ci_6144[4652];
	assign cj_6144[2933] = ci_6144[19];
	assign cj_6144[2934] = ci_6144[2490];
	assign cj_6144[2935] = ci_6144[5921];
	assign cj_6144[2936] = ci_6144[4168];
	assign cj_6144[2937] = ci_6144[3375];
	assign cj_6144[2938] = ci_6144[3542];
	assign cj_6144[2939] = ci_6144[4669];
	assign cj_6144[2940] = ci_6144[612];
	assign cj_6144[2941] = ci_6144[3659];
	assign cj_6144[2942] = ci_6144[1522];
	assign cj_6144[2943] = ci_6144[345];
	assign cj_6144[2944] = ci_6144[128];
	assign cj_6144[2945] = ci_6144[871];
	assign cj_6144[2946] = ci_6144[2574];
	assign cj_6144[2947] = ci_6144[5237];
	assign cj_6144[2948] = ci_6144[2716];
	assign cj_6144[2949] = ci_6144[1155];
	assign cj_6144[2950] = ci_6144[554];
	assign cj_6144[2951] = ci_6144[913];
	assign cj_6144[2952] = ci_6144[2232];
	assign cj_6144[2953] = ci_6144[4511];
	assign cj_6144[2954] = ci_6144[1606];
	assign cj_6144[2955] = ci_6144[5805];
	assign cj_6144[2956] = ci_6144[4820];
	assign cj_6144[2957] = ci_6144[4795];
	assign cj_6144[2958] = ci_6144[5730];
	assign cj_6144[2959] = ci_6144[1481];
	assign cj_6144[2960] = ci_6144[4336];
	assign cj_6144[2961] = ci_6144[2007];
	assign cj_6144[2962] = ci_6144[638];
	assign cj_6144[2963] = ci_6144[229];
	assign cj_6144[2964] = ci_6144[780];
	assign cj_6144[2965] = ci_6144[2291];
	assign cj_6144[2966] = ci_6144[4762];
	assign cj_6144[2967] = ci_6144[2049];
	assign cj_6144[2968] = ci_6144[296];
	assign cj_6144[2969] = ci_6144[5647];
	assign cj_6144[2970] = ci_6144[5814];
	assign cj_6144[2971] = ci_6144[797];
	assign cj_6144[2972] = ci_6144[2884];
	assign cj_6144[2973] = ci_6144[5931];
	assign cj_6144[2974] = ci_6144[3794];
	assign cj_6144[2975] = ci_6144[2617];
	assign cj_6144[2976] = ci_6144[2400];
	assign cj_6144[2977] = ci_6144[3143];
	assign cj_6144[2978] = ci_6144[4846];
	assign cj_6144[2979] = ci_6144[1365];
	assign cj_6144[2980] = ci_6144[4988];
	assign cj_6144[2981] = ci_6144[3427];
	assign cj_6144[2982] = ci_6144[2826];
	assign cj_6144[2983] = ci_6144[3185];
	assign cj_6144[2984] = ci_6144[4504];
	assign cj_6144[2985] = ci_6144[639];
	assign cj_6144[2986] = ci_6144[3878];
	assign cj_6144[2987] = ci_6144[1933];
	assign cj_6144[2988] = ci_6144[948];
	assign cj_6144[2989] = ci_6144[923];
	assign cj_6144[2990] = ci_6144[1858];
	assign cj_6144[2991] = ci_6144[3753];
	assign cj_6144[2992] = ci_6144[464];
	assign cj_6144[2993] = ci_6144[4279];
	assign cj_6144[2994] = ci_6144[2910];
	assign cj_6144[2995] = ci_6144[2501];
	assign cj_6144[2996] = ci_6144[3052];
	assign cj_6144[2997] = ci_6144[4563];
	assign cj_6144[2998] = ci_6144[890];
	assign cj_6144[2999] = ci_6144[4321];
	assign cj_6144[3000] = ci_6144[2568];
	assign cj_6144[3001] = ci_6144[1775];
	assign cj_6144[3002] = ci_6144[1942];
	assign cj_6144[3003] = ci_6144[3069];
	assign cj_6144[3004] = ci_6144[5156];
	assign cj_6144[3005] = ci_6144[2059];
	assign cj_6144[3006] = ci_6144[6066];
	assign cj_6144[3007] = ci_6144[4889];
	assign cj_6144[3008] = ci_6144[4672];
	assign cj_6144[3009] = ci_6144[5415];
	assign cj_6144[3010] = ci_6144[974];
	assign cj_6144[3011] = ci_6144[3637];
	assign cj_6144[3012] = ci_6144[1116];
	assign cj_6144[3013] = ci_6144[5699];
	assign cj_6144[3014] = ci_6144[5098];
	assign cj_6144[3015] = ci_6144[5457];
	assign cj_6144[3016] = ci_6144[632];
	assign cj_6144[3017] = ci_6144[2911];
	assign cj_6144[3018] = ci_6144[6];
	assign cj_6144[3019] = ci_6144[4205];
	assign cj_6144[3020] = ci_6144[3220];
	assign cj_6144[3021] = ci_6144[3195];
	assign cj_6144[3022] = ci_6144[4130];
	assign cj_6144[3023] = ci_6144[6025];
	assign cj_6144[3024] = ci_6144[2736];
	assign cj_6144[3025] = ci_6144[407];
	assign cj_6144[3026] = ci_6144[5182];
	assign cj_6144[3027] = ci_6144[4773];
	assign cj_6144[3028] = ci_6144[5324];
	assign cj_6144[3029] = ci_6144[691];
	assign cj_6144[3030] = ci_6144[3162];
	assign cj_6144[3031] = ci_6144[449];
	assign cj_6144[3032] = ci_6144[4840];
	assign cj_6144[3033] = ci_6144[4047];
	assign cj_6144[3034] = ci_6144[4214];
	assign cj_6144[3035] = ci_6144[5341];
	assign cj_6144[3036] = ci_6144[1284];
	assign cj_6144[3037] = ci_6144[4331];
	assign cj_6144[3038] = ci_6144[2194];
	assign cj_6144[3039] = ci_6144[1017];
	assign cj_6144[3040] = ci_6144[800];
	assign cj_6144[3041] = ci_6144[1543];
	assign cj_6144[3042] = ci_6144[3246];
	assign cj_6144[3043] = ci_6144[5909];
	assign cj_6144[3044] = ci_6144[3388];
	assign cj_6144[3045] = ci_6144[1827];
	assign cj_6144[3046] = ci_6144[1226];
	assign cj_6144[3047] = ci_6144[1585];
	assign cj_6144[3048] = ci_6144[2904];
	assign cj_6144[3049] = ci_6144[5183];
	assign cj_6144[3050] = ci_6144[2278];
	assign cj_6144[3051] = ci_6144[333];
	assign cj_6144[3052] = ci_6144[5492];
	assign cj_6144[3053] = ci_6144[5467];
	assign cj_6144[3054] = ci_6144[258];
	assign cj_6144[3055] = ci_6144[2153];
	assign cj_6144[3056] = ci_6144[5008];
	assign cj_6144[3057] = ci_6144[2679];
	assign cj_6144[3058] = ci_6144[1310];
	assign cj_6144[3059] = ci_6144[901];
	assign cj_6144[3060] = ci_6144[1452];
	assign cj_6144[3061] = ci_6144[2963];
	assign cj_6144[3062] = ci_6144[5434];
	assign cj_6144[3063] = ci_6144[2721];
	assign cj_6144[3064] = ci_6144[968];
	assign cj_6144[3065] = ci_6144[175];
	assign cj_6144[3066] = ci_6144[342];
	assign cj_6144[3067] = ci_6144[1469];
	assign cj_6144[3068] = ci_6144[3556];
	assign cj_6144[3069] = ci_6144[459];
	assign cj_6144[3070] = ci_6144[4466];
	assign cj_6144[3071] = ci_6144[3289];
	assign cj_6144[3072] = ci_6144[3072];
	assign cj_6144[3073] = ci_6144[3815];
	assign cj_6144[3074] = ci_6144[5518];
	assign cj_6144[3075] = ci_6144[2037];
	assign cj_6144[3076] = ci_6144[5660];
	assign cj_6144[3077] = ci_6144[4099];
	assign cj_6144[3078] = ci_6144[3498];
	assign cj_6144[3079] = ci_6144[3857];
	assign cj_6144[3080] = ci_6144[5176];
	assign cj_6144[3081] = ci_6144[1311];
	assign cj_6144[3082] = ci_6144[4550];
	assign cj_6144[3083] = ci_6144[2605];
	assign cj_6144[3084] = ci_6144[1620];
	assign cj_6144[3085] = ci_6144[1595];
	assign cj_6144[3086] = ci_6144[2530];
	assign cj_6144[3087] = ci_6144[4425];
	assign cj_6144[3088] = ci_6144[1136];
	assign cj_6144[3089] = ci_6144[4951];
	assign cj_6144[3090] = ci_6144[3582];
	assign cj_6144[3091] = ci_6144[3173];
	assign cj_6144[3092] = ci_6144[3724];
	assign cj_6144[3093] = ci_6144[5235];
	assign cj_6144[3094] = ci_6144[1562];
	assign cj_6144[3095] = ci_6144[4993];
	assign cj_6144[3096] = ci_6144[3240];
	assign cj_6144[3097] = ci_6144[2447];
	assign cj_6144[3098] = ci_6144[2614];
	assign cj_6144[3099] = ci_6144[3741];
	assign cj_6144[3100] = ci_6144[5828];
	assign cj_6144[3101] = ci_6144[2731];
	assign cj_6144[3102] = ci_6144[594];
	assign cj_6144[3103] = ci_6144[5561];
	assign cj_6144[3104] = ci_6144[5344];
	assign cj_6144[3105] = ci_6144[6087];
	assign cj_6144[3106] = ci_6144[1646];
	assign cj_6144[3107] = ci_6144[4309];
	assign cj_6144[3108] = ci_6144[1788];
	assign cj_6144[3109] = ci_6144[227];
	assign cj_6144[3110] = ci_6144[5770];
	assign cj_6144[3111] = ci_6144[6129];
	assign cj_6144[3112] = ci_6144[1304];
	assign cj_6144[3113] = ci_6144[3583];
	assign cj_6144[3114] = ci_6144[678];
	assign cj_6144[3115] = ci_6144[4877];
	assign cj_6144[3116] = ci_6144[3892];
	assign cj_6144[3117] = ci_6144[3867];
	assign cj_6144[3118] = ci_6144[4802];
	assign cj_6144[3119] = ci_6144[553];
	assign cj_6144[3120] = ci_6144[3408];
	assign cj_6144[3121] = ci_6144[1079];
	assign cj_6144[3122] = ci_6144[5854];
	assign cj_6144[3123] = ci_6144[5445];
	assign cj_6144[3124] = ci_6144[5996];
	assign cj_6144[3125] = ci_6144[1363];
	assign cj_6144[3126] = ci_6144[3834];
	assign cj_6144[3127] = ci_6144[1121];
	assign cj_6144[3128] = ci_6144[5512];
	assign cj_6144[3129] = ci_6144[4719];
	assign cj_6144[3130] = ci_6144[4886];
	assign cj_6144[3131] = ci_6144[6013];
	assign cj_6144[3132] = ci_6144[1956];
	assign cj_6144[3133] = ci_6144[5003];
	assign cj_6144[3134] = ci_6144[2866];
	assign cj_6144[3135] = ci_6144[1689];
	assign cj_6144[3136] = ci_6144[1472];
	assign cj_6144[3137] = ci_6144[2215];
	assign cj_6144[3138] = ci_6144[3918];
	assign cj_6144[3139] = ci_6144[437];
	assign cj_6144[3140] = ci_6144[4060];
	assign cj_6144[3141] = ci_6144[2499];
	assign cj_6144[3142] = ci_6144[1898];
	assign cj_6144[3143] = ci_6144[2257];
	assign cj_6144[3144] = ci_6144[3576];
	assign cj_6144[3145] = ci_6144[5855];
	assign cj_6144[3146] = ci_6144[2950];
	assign cj_6144[3147] = ci_6144[1005];
	assign cj_6144[3148] = ci_6144[20];
	assign cj_6144[3149] = ci_6144[6139];
	assign cj_6144[3150] = ci_6144[930];
	assign cj_6144[3151] = ci_6144[2825];
	assign cj_6144[3152] = ci_6144[5680];
	assign cj_6144[3153] = ci_6144[3351];
	assign cj_6144[3154] = ci_6144[1982];
	assign cj_6144[3155] = ci_6144[1573];
	assign cj_6144[3156] = ci_6144[2124];
	assign cj_6144[3157] = ci_6144[3635];
	assign cj_6144[3158] = ci_6144[6106];
	assign cj_6144[3159] = ci_6144[3393];
	assign cj_6144[3160] = ci_6144[1640];
	assign cj_6144[3161] = ci_6144[847];
	assign cj_6144[3162] = ci_6144[1014];
	assign cj_6144[3163] = ci_6144[2141];
	assign cj_6144[3164] = ci_6144[4228];
	assign cj_6144[3165] = ci_6144[1131];
	assign cj_6144[3166] = ci_6144[5138];
	assign cj_6144[3167] = ci_6144[3961];
	assign cj_6144[3168] = ci_6144[3744];
	assign cj_6144[3169] = ci_6144[4487];
	assign cj_6144[3170] = ci_6144[46];
	assign cj_6144[3171] = ci_6144[2709];
	assign cj_6144[3172] = ci_6144[188];
	assign cj_6144[3173] = ci_6144[4771];
	assign cj_6144[3174] = ci_6144[4170];
	assign cj_6144[3175] = ci_6144[4529];
	assign cj_6144[3176] = ci_6144[5848];
	assign cj_6144[3177] = ci_6144[1983];
	assign cj_6144[3178] = ci_6144[5222];
	assign cj_6144[3179] = ci_6144[3277];
	assign cj_6144[3180] = ci_6144[2292];
	assign cj_6144[3181] = ci_6144[2267];
	assign cj_6144[3182] = ci_6144[3202];
	assign cj_6144[3183] = ci_6144[5097];
	assign cj_6144[3184] = ci_6144[1808];
	assign cj_6144[3185] = ci_6144[5623];
	assign cj_6144[3186] = ci_6144[4254];
	assign cj_6144[3187] = ci_6144[3845];
	assign cj_6144[3188] = ci_6144[4396];
	assign cj_6144[3189] = ci_6144[5907];
	assign cj_6144[3190] = ci_6144[2234];
	assign cj_6144[3191] = ci_6144[5665];
	assign cj_6144[3192] = ci_6144[3912];
	assign cj_6144[3193] = ci_6144[3119];
	assign cj_6144[3194] = ci_6144[3286];
	assign cj_6144[3195] = ci_6144[4413];
	assign cj_6144[3196] = ci_6144[356];
	assign cj_6144[3197] = ci_6144[3403];
	assign cj_6144[3198] = ci_6144[1266];
	assign cj_6144[3199] = ci_6144[89];
	assign cj_6144[3200] = ci_6144[6016];
	assign cj_6144[3201] = ci_6144[615];
	assign cj_6144[3202] = ci_6144[2318];
	assign cj_6144[3203] = ci_6144[4981];
	assign cj_6144[3204] = ci_6144[2460];
	assign cj_6144[3205] = ci_6144[899];
	assign cj_6144[3206] = ci_6144[298];
	assign cj_6144[3207] = ci_6144[657];
	assign cj_6144[3208] = ci_6144[1976];
	assign cj_6144[3209] = ci_6144[4255];
	assign cj_6144[3210] = ci_6144[1350];
	assign cj_6144[3211] = ci_6144[5549];
	assign cj_6144[3212] = ci_6144[4564];
	assign cj_6144[3213] = ci_6144[4539];
	assign cj_6144[3214] = ci_6144[5474];
	assign cj_6144[3215] = ci_6144[1225];
	assign cj_6144[3216] = ci_6144[4080];
	assign cj_6144[3217] = ci_6144[1751];
	assign cj_6144[3218] = ci_6144[382];
	assign cj_6144[3219] = ci_6144[6117];
	assign cj_6144[3220] = ci_6144[524];
	assign cj_6144[3221] = ci_6144[2035];
	assign cj_6144[3222] = ci_6144[4506];
	assign cj_6144[3223] = ci_6144[1793];
	assign cj_6144[3224] = ci_6144[40];
	assign cj_6144[3225] = ci_6144[5391];
	assign cj_6144[3226] = ci_6144[5558];
	assign cj_6144[3227] = ci_6144[541];
	assign cj_6144[3228] = ci_6144[2628];
	assign cj_6144[3229] = ci_6144[5675];
	assign cj_6144[3230] = ci_6144[3538];
	assign cj_6144[3231] = ci_6144[2361];
	assign cj_6144[3232] = ci_6144[2144];
	assign cj_6144[3233] = ci_6144[2887];
	assign cj_6144[3234] = ci_6144[4590];
	assign cj_6144[3235] = ci_6144[1109];
	assign cj_6144[3236] = ci_6144[4732];
	assign cj_6144[3237] = ci_6144[3171];
	assign cj_6144[3238] = ci_6144[2570];
	assign cj_6144[3239] = ci_6144[2929];
	assign cj_6144[3240] = ci_6144[4248];
	assign cj_6144[3241] = ci_6144[383];
	assign cj_6144[3242] = ci_6144[3622];
	assign cj_6144[3243] = ci_6144[1677];
	assign cj_6144[3244] = ci_6144[692];
	assign cj_6144[3245] = ci_6144[667];
	assign cj_6144[3246] = ci_6144[1602];
	assign cj_6144[3247] = ci_6144[3497];
	assign cj_6144[3248] = ci_6144[208];
	assign cj_6144[3249] = ci_6144[4023];
	assign cj_6144[3250] = ci_6144[2654];
	assign cj_6144[3251] = ci_6144[2245];
	assign cj_6144[3252] = ci_6144[2796];
	assign cj_6144[3253] = ci_6144[4307];
	assign cj_6144[3254] = ci_6144[634];
	assign cj_6144[3255] = ci_6144[4065];
	assign cj_6144[3256] = ci_6144[2312];
	assign cj_6144[3257] = ci_6144[1519];
	assign cj_6144[3258] = ci_6144[1686];
	assign cj_6144[3259] = ci_6144[2813];
	assign cj_6144[3260] = ci_6144[4900];
	assign cj_6144[3261] = ci_6144[1803];
	assign cj_6144[3262] = ci_6144[5810];
	assign cj_6144[3263] = ci_6144[4633];
	assign cj_6144[3264] = ci_6144[4416];
	assign cj_6144[3265] = ci_6144[5159];
	assign cj_6144[3266] = ci_6144[718];
	assign cj_6144[3267] = ci_6144[3381];
	assign cj_6144[3268] = ci_6144[860];
	assign cj_6144[3269] = ci_6144[5443];
	assign cj_6144[3270] = ci_6144[4842];
	assign cj_6144[3271] = ci_6144[5201];
	assign cj_6144[3272] = ci_6144[376];
	assign cj_6144[3273] = ci_6144[2655];
	assign cj_6144[3274] = ci_6144[5894];
	assign cj_6144[3275] = ci_6144[3949];
	assign cj_6144[3276] = ci_6144[2964];
	assign cj_6144[3277] = ci_6144[2939];
	assign cj_6144[3278] = ci_6144[3874];
	assign cj_6144[3279] = ci_6144[5769];
	assign cj_6144[3280] = ci_6144[2480];
	assign cj_6144[3281] = ci_6144[151];
	assign cj_6144[3282] = ci_6144[4926];
	assign cj_6144[3283] = ci_6144[4517];
	assign cj_6144[3284] = ci_6144[5068];
	assign cj_6144[3285] = ci_6144[435];
	assign cj_6144[3286] = ci_6144[2906];
	assign cj_6144[3287] = ci_6144[193];
	assign cj_6144[3288] = ci_6144[4584];
	assign cj_6144[3289] = ci_6144[3791];
	assign cj_6144[3290] = ci_6144[3958];
	assign cj_6144[3291] = ci_6144[5085];
	assign cj_6144[3292] = ci_6144[1028];
	assign cj_6144[3293] = ci_6144[4075];
	assign cj_6144[3294] = ci_6144[1938];
	assign cj_6144[3295] = ci_6144[761];
	assign cj_6144[3296] = ci_6144[544];
	assign cj_6144[3297] = ci_6144[1287];
	assign cj_6144[3298] = ci_6144[2990];
	assign cj_6144[3299] = ci_6144[5653];
	assign cj_6144[3300] = ci_6144[3132];
	assign cj_6144[3301] = ci_6144[1571];
	assign cj_6144[3302] = ci_6144[970];
	assign cj_6144[3303] = ci_6144[1329];
	assign cj_6144[3304] = ci_6144[2648];
	assign cj_6144[3305] = ci_6144[4927];
	assign cj_6144[3306] = ci_6144[2022];
	assign cj_6144[3307] = ci_6144[77];
	assign cj_6144[3308] = ci_6144[5236];
	assign cj_6144[3309] = ci_6144[5211];
	assign cj_6144[3310] = ci_6144[2];
	assign cj_6144[3311] = ci_6144[1897];
	assign cj_6144[3312] = ci_6144[4752];
	assign cj_6144[3313] = ci_6144[2423];
	assign cj_6144[3314] = ci_6144[1054];
	assign cj_6144[3315] = ci_6144[645];
	assign cj_6144[3316] = ci_6144[1196];
	assign cj_6144[3317] = ci_6144[2707];
	assign cj_6144[3318] = ci_6144[5178];
	assign cj_6144[3319] = ci_6144[2465];
	assign cj_6144[3320] = ci_6144[712];
	assign cj_6144[3321] = ci_6144[6063];
	assign cj_6144[3322] = ci_6144[86];
	assign cj_6144[3323] = ci_6144[1213];
	assign cj_6144[3324] = ci_6144[3300];
	assign cj_6144[3325] = ci_6144[203];
	assign cj_6144[3326] = ci_6144[4210];
	assign cj_6144[3327] = ci_6144[3033];
	assign cj_6144[3328] = ci_6144[2816];
	assign cj_6144[3329] = ci_6144[3559];
	assign cj_6144[3330] = ci_6144[5262];
	assign cj_6144[3331] = ci_6144[1781];
	assign cj_6144[3332] = ci_6144[5404];
	assign cj_6144[3333] = ci_6144[3843];
	assign cj_6144[3334] = ci_6144[3242];
	assign cj_6144[3335] = ci_6144[3601];
	assign cj_6144[3336] = ci_6144[4920];
	assign cj_6144[3337] = ci_6144[1055];
	assign cj_6144[3338] = ci_6144[4294];
	assign cj_6144[3339] = ci_6144[2349];
	assign cj_6144[3340] = ci_6144[1364];
	assign cj_6144[3341] = ci_6144[1339];
	assign cj_6144[3342] = ci_6144[2274];
	assign cj_6144[3343] = ci_6144[4169];
	assign cj_6144[3344] = ci_6144[880];
	assign cj_6144[3345] = ci_6144[4695];
	assign cj_6144[3346] = ci_6144[3326];
	assign cj_6144[3347] = ci_6144[2917];
	assign cj_6144[3348] = ci_6144[3468];
	assign cj_6144[3349] = ci_6144[4979];
	assign cj_6144[3350] = ci_6144[1306];
	assign cj_6144[3351] = ci_6144[4737];
	assign cj_6144[3352] = ci_6144[2984];
	assign cj_6144[3353] = ci_6144[2191];
	assign cj_6144[3354] = ci_6144[2358];
	assign cj_6144[3355] = ci_6144[3485];
	assign cj_6144[3356] = ci_6144[5572];
	assign cj_6144[3357] = ci_6144[2475];
	assign cj_6144[3358] = ci_6144[338];
	assign cj_6144[3359] = ci_6144[5305];
	assign cj_6144[3360] = ci_6144[5088];
	assign cj_6144[3361] = ci_6144[5831];
	assign cj_6144[3362] = ci_6144[1390];
	assign cj_6144[3363] = ci_6144[4053];
	assign cj_6144[3364] = ci_6144[1532];
	assign cj_6144[3365] = ci_6144[6115];
	assign cj_6144[3366] = ci_6144[5514];
	assign cj_6144[3367] = ci_6144[5873];
	assign cj_6144[3368] = ci_6144[1048];
	assign cj_6144[3369] = ci_6144[3327];
	assign cj_6144[3370] = ci_6144[422];
	assign cj_6144[3371] = ci_6144[4621];
	assign cj_6144[3372] = ci_6144[3636];
	assign cj_6144[3373] = ci_6144[3611];
	assign cj_6144[3374] = ci_6144[4546];
	assign cj_6144[3375] = ci_6144[297];
	assign cj_6144[3376] = ci_6144[3152];
	assign cj_6144[3377] = ci_6144[823];
	assign cj_6144[3378] = ci_6144[5598];
	assign cj_6144[3379] = ci_6144[5189];
	assign cj_6144[3380] = ci_6144[5740];
	assign cj_6144[3381] = ci_6144[1107];
	assign cj_6144[3382] = ci_6144[3578];
	assign cj_6144[3383] = ci_6144[865];
	assign cj_6144[3384] = ci_6144[5256];
	assign cj_6144[3385] = ci_6144[4463];
	assign cj_6144[3386] = ci_6144[4630];
	assign cj_6144[3387] = ci_6144[5757];
	assign cj_6144[3388] = ci_6144[1700];
	assign cj_6144[3389] = ci_6144[4747];
	assign cj_6144[3390] = ci_6144[2610];
	assign cj_6144[3391] = ci_6144[1433];
	assign cj_6144[3392] = ci_6144[1216];
	assign cj_6144[3393] = ci_6144[1959];
	assign cj_6144[3394] = ci_6144[3662];
	assign cj_6144[3395] = ci_6144[181];
	assign cj_6144[3396] = ci_6144[3804];
	assign cj_6144[3397] = ci_6144[2243];
	assign cj_6144[3398] = ci_6144[1642];
	assign cj_6144[3399] = ci_6144[2001];
	assign cj_6144[3400] = ci_6144[3320];
	assign cj_6144[3401] = ci_6144[5599];
	assign cj_6144[3402] = ci_6144[2694];
	assign cj_6144[3403] = ci_6144[749];
	assign cj_6144[3404] = ci_6144[5908];
	assign cj_6144[3405] = ci_6144[5883];
	assign cj_6144[3406] = ci_6144[674];
	assign cj_6144[3407] = ci_6144[2569];
	assign cj_6144[3408] = ci_6144[5424];
	assign cj_6144[3409] = ci_6144[3095];
	assign cj_6144[3410] = ci_6144[1726];
	assign cj_6144[3411] = ci_6144[1317];
	assign cj_6144[3412] = ci_6144[1868];
	assign cj_6144[3413] = ci_6144[3379];
	assign cj_6144[3414] = ci_6144[5850];
	assign cj_6144[3415] = ci_6144[3137];
	assign cj_6144[3416] = ci_6144[1384];
	assign cj_6144[3417] = ci_6144[591];
	assign cj_6144[3418] = ci_6144[758];
	assign cj_6144[3419] = ci_6144[1885];
	assign cj_6144[3420] = ci_6144[3972];
	assign cj_6144[3421] = ci_6144[875];
	assign cj_6144[3422] = ci_6144[4882];
	assign cj_6144[3423] = ci_6144[3705];
	assign cj_6144[3424] = ci_6144[3488];
	assign cj_6144[3425] = ci_6144[4231];
	assign cj_6144[3426] = ci_6144[5934];
	assign cj_6144[3427] = ci_6144[2453];
	assign cj_6144[3428] = ci_6144[6076];
	assign cj_6144[3429] = ci_6144[4515];
	assign cj_6144[3430] = ci_6144[3914];
	assign cj_6144[3431] = ci_6144[4273];
	assign cj_6144[3432] = ci_6144[5592];
	assign cj_6144[3433] = ci_6144[1727];
	assign cj_6144[3434] = ci_6144[4966];
	assign cj_6144[3435] = ci_6144[3021];
	assign cj_6144[3436] = ci_6144[2036];
	assign cj_6144[3437] = ci_6144[2011];
	assign cj_6144[3438] = ci_6144[2946];
	assign cj_6144[3439] = ci_6144[4841];
	assign cj_6144[3440] = ci_6144[1552];
	assign cj_6144[3441] = ci_6144[5367];
	assign cj_6144[3442] = ci_6144[3998];
	assign cj_6144[3443] = ci_6144[3589];
	assign cj_6144[3444] = ci_6144[4140];
	assign cj_6144[3445] = ci_6144[5651];
	assign cj_6144[3446] = ci_6144[1978];
	assign cj_6144[3447] = ci_6144[5409];
	assign cj_6144[3448] = ci_6144[3656];
	assign cj_6144[3449] = ci_6144[2863];
	assign cj_6144[3450] = ci_6144[3030];
	assign cj_6144[3451] = ci_6144[4157];
	assign cj_6144[3452] = ci_6144[100];
	assign cj_6144[3453] = ci_6144[3147];
	assign cj_6144[3454] = ci_6144[1010];
	assign cj_6144[3455] = ci_6144[5977];
	assign cj_6144[3456] = ci_6144[5760];
	assign cj_6144[3457] = ci_6144[359];
	assign cj_6144[3458] = ci_6144[2062];
	assign cj_6144[3459] = ci_6144[4725];
	assign cj_6144[3460] = ci_6144[2204];
	assign cj_6144[3461] = ci_6144[643];
	assign cj_6144[3462] = ci_6144[42];
	assign cj_6144[3463] = ci_6144[401];
	assign cj_6144[3464] = ci_6144[1720];
	assign cj_6144[3465] = ci_6144[3999];
	assign cj_6144[3466] = ci_6144[1094];
	assign cj_6144[3467] = ci_6144[5293];
	assign cj_6144[3468] = ci_6144[4308];
	assign cj_6144[3469] = ci_6144[4283];
	assign cj_6144[3470] = ci_6144[5218];
	assign cj_6144[3471] = ci_6144[969];
	assign cj_6144[3472] = ci_6144[3824];
	assign cj_6144[3473] = ci_6144[1495];
	assign cj_6144[3474] = ci_6144[126];
	assign cj_6144[3475] = ci_6144[5861];
	assign cj_6144[3476] = ci_6144[268];
	assign cj_6144[3477] = ci_6144[1779];
	assign cj_6144[3478] = ci_6144[4250];
	assign cj_6144[3479] = ci_6144[1537];
	assign cj_6144[3480] = ci_6144[5928];
	assign cj_6144[3481] = ci_6144[5135];
	assign cj_6144[3482] = ci_6144[5302];
	assign cj_6144[3483] = ci_6144[285];
	assign cj_6144[3484] = ci_6144[2372];
	assign cj_6144[3485] = ci_6144[5419];
	assign cj_6144[3486] = ci_6144[3282];
	assign cj_6144[3487] = ci_6144[2105];
	assign cj_6144[3488] = ci_6144[1888];
	assign cj_6144[3489] = ci_6144[2631];
	assign cj_6144[3490] = ci_6144[4334];
	assign cj_6144[3491] = ci_6144[853];
	assign cj_6144[3492] = ci_6144[4476];
	assign cj_6144[3493] = ci_6144[2915];
	assign cj_6144[3494] = ci_6144[2314];
	assign cj_6144[3495] = ci_6144[2673];
	assign cj_6144[3496] = ci_6144[3992];
	assign cj_6144[3497] = ci_6144[127];
	assign cj_6144[3498] = ci_6144[3366];
	assign cj_6144[3499] = ci_6144[1421];
	assign cj_6144[3500] = ci_6144[436];
	assign cj_6144[3501] = ci_6144[411];
	assign cj_6144[3502] = ci_6144[1346];
	assign cj_6144[3503] = ci_6144[3241];
	assign cj_6144[3504] = ci_6144[6096];
	assign cj_6144[3505] = ci_6144[3767];
	assign cj_6144[3506] = ci_6144[2398];
	assign cj_6144[3507] = ci_6144[1989];
	assign cj_6144[3508] = ci_6144[2540];
	assign cj_6144[3509] = ci_6144[4051];
	assign cj_6144[3510] = ci_6144[378];
	assign cj_6144[3511] = ci_6144[3809];
	assign cj_6144[3512] = ci_6144[2056];
	assign cj_6144[3513] = ci_6144[1263];
	assign cj_6144[3514] = ci_6144[1430];
	assign cj_6144[3515] = ci_6144[2557];
	assign cj_6144[3516] = ci_6144[4644];
	assign cj_6144[3517] = ci_6144[1547];
	assign cj_6144[3518] = ci_6144[5554];
	assign cj_6144[3519] = ci_6144[4377];
	assign cj_6144[3520] = ci_6144[4160];
	assign cj_6144[3521] = ci_6144[4903];
	assign cj_6144[3522] = ci_6144[462];
	assign cj_6144[3523] = ci_6144[3125];
	assign cj_6144[3524] = ci_6144[604];
	assign cj_6144[3525] = ci_6144[5187];
	assign cj_6144[3526] = ci_6144[4586];
	assign cj_6144[3527] = ci_6144[4945];
	assign cj_6144[3528] = ci_6144[120];
	assign cj_6144[3529] = ci_6144[2399];
	assign cj_6144[3530] = ci_6144[5638];
	assign cj_6144[3531] = ci_6144[3693];
	assign cj_6144[3532] = ci_6144[2708];
	assign cj_6144[3533] = ci_6144[2683];
	assign cj_6144[3534] = ci_6144[3618];
	assign cj_6144[3535] = ci_6144[5513];
	assign cj_6144[3536] = ci_6144[2224];
	assign cj_6144[3537] = ci_6144[6039];
	assign cj_6144[3538] = ci_6144[4670];
	assign cj_6144[3539] = ci_6144[4261];
	assign cj_6144[3540] = ci_6144[4812];
	assign cj_6144[3541] = ci_6144[179];
	assign cj_6144[3542] = ci_6144[2650];
	assign cj_6144[3543] = ci_6144[6081];
	assign cj_6144[3544] = ci_6144[4328];
	assign cj_6144[3545] = ci_6144[3535];
	assign cj_6144[3546] = ci_6144[3702];
	assign cj_6144[3547] = ci_6144[4829];
	assign cj_6144[3548] = ci_6144[772];
	assign cj_6144[3549] = ci_6144[3819];
	assign cj_6144[3550] = ci_6144[1682];
	assign cj_6144[3551] = ci_6144[505];
	assign cj_6144[3552] = ci_6144[288];
	assign cj_6144[3553] = ci_6144[1031];
	assign cj_6144[3554] = ci_6144[2734];
	assign cj_6144[3555] = ci_6144[5397];
	assign cj_6144[3556] = ci_6144[2876];
	assign cj_6144[3557] = ci_6144[1315];
	assign cj_6144[3558] = ci_6144[714];
	assign cj_6144[3559] = ci_6144[1073];
	assign cj_6144[3560] = ci_6144[2392];
	assign cj_6144[3561] = ci_6144[4671];
	assign cj_6144[3562] = ci_6144[1766];
	assign cj_6144[3563] = ci_6144[5965];
	assign cj_6144[3564] = ci_6144[4980];
	assign cj_6144[3565] = ci_6144[4955];
	assign cj_6144[3566] = ci_6144[5890];
	assign cj_6144[3567] = ci_6144[1641];
	assign cj_6144[3568] = ci_6144[4496];
	assign cj_6144[3569] = ci_6144[2167];
	assign cj_6144[3570] = ci_6144[798];
	assign cj_6144[3571] = ci_6144[389];
	assign cj_6144[3572] = ci_6144[940];
	assign cj_6144[3573] = ci_6144[2451];
	assign cj_6144[3574] = ci_6144[4922];
	assign cj_6144[3575] = ci_6144[2209];
	assign cj_6144[3576] = ci_6144[456];
	assign cj_6144[3577] = ci_6144[5807];
	assign cj_6144[3578] = ci_6144[5974];
	assign cj_6144[3579] = ci_6144[957];
	assign cj_6144[3580] = ci_6144[3044];
	assign cj_6144[3581] = ci_6144[6091];
	assign cj_6144[3582] = ci_6144[3954];
	assign cj_6144[3583] = ci_6144[2777];
	assign cj_6144[3584] = ci_6144[2560];
	assign cj_6144[3585] = ci_6144[3303];
	assign cj_6144[3586] = ci_6144[5006];
	assign cj_6144[3587] = ci_6144[1525];
	assign cj_6144[3588] = ci_6144[5148];
	assign cj_6144[3589] = ci_6144[3587];
	assign cj_6144[3590] = ci_6144[2986];
	assign cj_6144[3591] = ci_6144[3345];
	assign cj_6144[3592] = ci_6144[4664];
	assign cj_6144[3593] = ci_6144[799];
	assign cj_6144[3594] = ci_6144[4038];
	assign cj_6144[3595] = ci_6144[2093];
	assign cj_6144[3596] = ci_6144[1108];
	assign cj_6144[3597] = ci_6144[1083];
	assign cj_6144[3598] = ci_6144[2018];
	assign cj_6144[3599] = ci_6144[3913];
	assign cj_6144[3600] = ci_6144[624];
	assign cj_6144[3601] = ci_6144[4439];
	assign cj_6144[3602] = ci_6144[3070];
	assign cj_6144[3603] = ci_6144[2661];
	assign cj_6144[3604] = ci_6144[3212];
	assign cj_6144[3605] = ci_6144[4723];
	assign cj_6144[3606] = ci_6144[1050];
	assign cj_6144[3607] = ci_6144[4481];
	assign cj_6144[3608] = ci_6144[2728];
	assign cj_6144[3609] = ci_6144[1935];
	assign cj_6144[3610] = ci_6144[2102];
	assign cj_6144[3611] = ci_6144[3229];
	assign cj_6144[3612] = ci_6144[5316];
	assign cj_6144[3613] = ci_6144[2219];
	assign cj_6144[3614] = ci_6144[82];
	assign cj_6144[3615] = ci_6144[5049];
	assign cj_6144[3616] = ci_6144[4832];
	assign cj_6144[3617] = ci_6144[5575];
	assign cj_6144[3618] = ci_6144[1134];
	assign cj_6144[3619] = ci_6144[3797];
	assign cj_6144[3620] = ci_6144[1276];
	assign cj_6144[3621] = ci_6144[5859];
	assign cj_6144[3622] = ci_6144[5258];
	assign cj_6144[3623] = ci_6144[5617];
	assign cj_6144[3624] = ci_6144[792];
	assign cj_6144[3625] = ci_6144[3071];
	assign cj_6144[3626] = ci_6144[166];
	assign cj_6144[3627] = ci_6144[4365];
	assign cj_6144[3628] = ci_6144[3380];
	assign cj_6144[3629] = ci_6144[3355];
	assign cj_6144[3630] = ci_6144[4290];
	assign cj_6144[3631] = ci_6144[41];
	assign cj_6144[3632] = ci_6144[2896];
	assign cj_6144[3633] = ci_6144[567];
	assign cj_6144[3634] = ci_6144[5342];
	assign cj_6144[3635] = ci_6144[4933];
	assign cj_6144[3636] = ci_6144[5484];
	assign cj_6144[3637] = ci_6144[851];
	assign cj_6144[3638] = ci_6144[3322];
	assign cj_6144[3639] = ci_6144[609];
	assign cj_6144[3640] = ci_6144[5000];
	assign cj_6144[3641] = ci_6144[4207];
	assign cj_6144[3642] = ci_6144[4374];
	assign cj_6144[3643] = ci_6144[5501];
	assign cj_6144[3644] = ci_6144[1444];
	assign cj_6144[3645] = ci_6144[4491];
	assign cj_6144[3646] = ci_6144[2354];
	assign cj_6144[3647] = ci_6144[1177];
	assign cj_6144[3648] = ci_6144[960];
	assign cj_6144[3649] = ci_6144[1703];
	assign cj_6144[3650] = ci_6144[3406];
	assign cj_6144[3651] = ci_6144[6069];
	assign cj_6144[3652] = ci_6144[3548];
	assign cj_6144[3653] = ci_6144[1987];
	assign cj_6144[3654] = ci_6144[1386];
	assign cj_6144[3655] = ci_6144[1745];
	assign cj_6144[3656] = ci_6144[3064];
	assign cj_6144[3657] = ci_6144[5343];
	assign cj_6144[3658] = ci_6144[2438];
	assign cj_6144[3659] = ci_6144[493];
	assign cj_6144[3660] = ci_6144[5652];
	assign cj_6144[3661] = ci_6144[5627];
	assign cj_6144[3662] = ci_6144[418];
	assign cj_6144[3663] = ci_6144[2313];
	assign cj_6144[3664] = ci_6144[5168];
	assign cj_6144[3665] = ci_6144[2839];
	assign cj_6144[3666] = ci_6144[1470];
	assign cj_6144[3667] = ci_6144[1061];
	assign cj_6144[3668] = ci_6144[1612];
	assign cj_6144[3669] = ci_6144[3123];
	assign cj_6144[3670] = ci_6144[5594];
	assign cj_6144[3671] = ci_6144[2881];
	assign cj_6144[3672] = ci_6144[1128];
	assign cj_6144[3673] = ci_6144[335];
	assign cj_6144[3674] = ci_6144[502];
	assign cj_6144[3675] = ci_6144[1629];
	assign cj_6144[3676] = ci_6144[3716];
	assign cj_6144[3677] = ci_6144[619];
	assign cj_6144[3678] = ci_6144[4626];
	assign cj_6144[3679] = ci_6144[3449];
	assign cj_6144[3680] = ci_6144[3232];
	assign cj_6144[3681] = ci_6144[3975];
	assign cj_6144[3682] = ci_6144[5678];
	assign cj_6144[3683] = ci_6144[2197];
	assign cj_6144[3684] = ci_6144[5820];
	assign cj_6144[3685] = ci_6144[4259];
	assign cj_6144[3686] = ci_6144[3658];
	assign cj_6144[3687] = ci_6144[4017];
	assign cj_6144[3688] = ci_6144[5336];
	assign cj_6144[3689] = ci_6144[1471];
	assign cj_6144[3690] = ci_6144[4710];
	assign cj_6144[3691] = ci_6144[2765];
	assign cj_6144[3692] = ci_6144[1780];
	assign cj_6144[3693] = ci_6144[1755];
	assign cj_6144[3694] = ci_6144[2690];
	assign cj_6144[3695] = ci_6144[4585];
	assign cj_6144[3696] = ci_6144[1296];
	assign cj_6144[3697] = ci_6144[5111];
	assign cj_6144[3698] = ci_6144[3742];
	assign cj_6144[3699] = ci_6144[3333];
	assign cj_6144[3700] = ci_6144[3884];
	assign cj_6144[3701] = ci_6144[5395];
	assign cj_6144[3702] = ci_6144[1722];
	assign cj_6144[3703] = ci_6144[5153];
	assign cj_6144[3704] = ci_6144[3400];
	assign cj_6144[3705] = ci_6144[2607];
	assign cj_6144[3706] = ci_6144[2774];
	assign cj_6144[3707] = ci_6144[3901];
	assign cj_6144[3708] = ci_6144[5988];
	assign cj_6144[3709] = ci_6144[2891];
	assign cj_6144[3710] = ci_6144[754];
	assign cj_6144[3711] = ci_6144[5721];
	assign cj_6144[3712] = ci_6144[5504];
	assign cj_6144[3713] = ci_6144[103];
	assign cj_6144[3714] = ci_6144[1806];
	assign cj_6144[3715] = ci_6144[4469];
	assign cj_6144[3716] = ci_6144[1948];
	assign cj_6144[3717] = ci_6144[387];
	assign cj_6144[3718] = ci_6144[5930];
	assign cj_6144[3719] = ci_6144[145];
	assign cj_6144[3720] = ci_6144[1464];
	assign cj_6144[3721] = ci_6144[3743];
	assign cj_6144[3722] = ci_6144[838];
	assign cj_6144[3723] = ci_6144[5037];
	assign cj_6144[3724] = ci_6144[4052];
	assign cj_6144[3725] = ci_6144[4027];
	assign cj_6144[3726] = ci_6144[4962];
	assign cj_6144[3727] = ci_6144[713];
	assign cj_6144[3728] = ci_6144[3568];
	assign cj_6144[3729] = ci_6144[1239];
	assign cj_6144[3730] = ci_6144[6014];
	assign cj_6144[3731] = ci_6144[5605];
	assign cj_6144[3732] = ci_6144[12];
	assign cj_6144[3733] = ci_6144[1523];
	assign cj_6144[3734] = ci_6144[3994];
	assign cj_6144[3735] = ci_6144[1281];
	assign cj_6144[3736] = ci_6144[5672];
	assign cj_6144[3737] = ci_6144[4879];
	assign cj_6144[3738] = ci_6144[5046];
	assign cj_6144[3739] = ci_6144[29];
	assign cj_6144[3740] = ci_6144[2116];
	assign cj_6144[3741] = ci_6144[5163];
	assign cj_6144[3742] = ci_6144[3026];
	assign cj_6144[3743] = ci_6144[1849];
	assign cj_6144[3744] = ci_6144[1632];
	assign cj_6144[3745] = ci_6144[2375];
	assign cj_6144[3746] = ci_6144[4078];
	assign cj_6144[3747] = ci_6144[597];
	assign cj_6144[3748] = ci_6144[4220];
	assign cj_6144[3749] = ci_6144[2659];
	assign cj_6144[3750] = ci_6144[2058];
	assign cj_6144[3751] = ci_6144[2417];
	assign cj_6144[3752] = ci_6144[3736];
	assign cj_6144[3753] = ci_6144[6015];
	assign cj_6144[3754] = ci_6144[3110];
	assign cj_6144[3755] = ci_6144[1165];
	assign cj_6144[3756] = ci_6144[180];
	assign cj_6144[3757] = ci_6144[155];
	assign cj_6144[3758] = ci_6144[1090];
	assign cj_6144[3759] = ci_6144[2985];
	assign cj_6144[3760] = ci_6144[5840];
	assign cj_6144[3761] = ci_6144[3511];
	assign cj_6144[3762] = ci_6144[2142];
	assign cj_6144[3763] = ci_6144[1733];
	assign cj_6144[3764] = ci_6144[2284];
	assign cj_6144[3765] = ci_6144[3795];
	assign cj_6144[3766] = ci_6144[122];
	assign cj_6144[3767] = ci_6144[3553];
	assign cj_6144[3768] = ci_6144[1800];
	assign cj_6144[3769] = ci_6144[1007];
	assign cj_6144[3770] = ci_6144[1174];
	assign cj_6144[3771] = ci_6144[2301];
	assign cj_6144[3772] = ci_6144[4388];
	assign cj_6144[3773] = ci_6144[1291];
	assign cj_6144[3774] = ci_6144[5298];
	assign cj_6144[3775] = ci_6144[4121];
	assign cj_6144[3776] = ci_6144[3904];
	assign cj_6144[3777] = ci_6144[4647];
	assign cj_6144[3778] = ci_6144[206];
	assign cj_6144[3779] = ci_6144[2869];
	assign cj_6144[3780] = ci_6144[348];
	assign cj_6144[3781] = ci_6144[4931];
	assign cj_6144[3782] = ci_6144[4330];
	assign cj_6144[3783] = ci_6144[4689];
	assign cj_6144[3784] = ci_6144[6008];
	assign cj_6144[3785] = ci_6144[2143];
	assign cj_6144[3786] = ci_6144[5382];
	assign cj_6144[3787] = ci_6144[3437];
	assign cj_6144[3788] = ci_6144[2452];
	assign cj_6144[3789] = ci_6144[2427];
	assign cj_6144[3790] = ci_6144[3362];
	assign cj_6144[3791] = ci_6144[5257];
	assign cj_6144[3792] = ci_6144[1968];
	assign cj_6144[3793] = ci_6144[5783];
	assign cj_6144[3794] = ci_6144[4414];
	assign cj_6144[3795] = ci_6144[4005];
	assign cj_6144[3796] = ci_6144[4556];
	assign cj_6144[3797] = ci_6144[6067];
	assign cj_6144[3798] = ci_6144[2394];
	assign cj_6144[3799] = ci_6144[5825];
	assign cj_6144[3800] = ci_6144[4072];
	assign cj_6144[3801] = ci_6144[3279];
	assign cj_6144[3802] = ci_6144[3446];
	assign cj_6144[3803] = ci_6144[4573];
	assign cj_6144[3804] = ci_6144[516];
	assign cj_6144[3805] = ci_6144[3563];
	assign cj_6144[3806] = ci_6144[1426];
	assign cj_6144[3807] = ci_6144[249];
	assign cj_6144[3808] = ci_6144[32];
	assign cj_6144[3809] = ci_6144[775];
	assign cj_6144[3810] = ci_6144[2478];
	assign cj_6144[3811] = ci_6144[5141];
	assign cj_6144[3812] = ci_6144[2620];
	assign cj_6144[3813] = ci_6144[1059];
	assign cj_6144[3814] = ci_6144[458];
	assign cj_6144[3815] = ci_6144[817];
	assign cj_6144[3816] = ci_6144[2136];
	assign cj_6144[3817] = ci_6144[4415];
	assign cj_6144[3818] = ci_6144[1510];
	assign cj_6144[3819] = ci_6144[5709];
	assign cj_6144[3820] = ci_6144[4724];
	assign cj_6144[3821] = ci_6144[4699];
	assign cj_6144[3822] = ci_6144[5634];
	assign cj_6144[3823] = ci_6144[1385];
	assign cj_6144[3824] = ci_6144[4240];
	assign cj_6144[3825] = ci_6144[1911];
	assign cj_6144[3826] = ci_6144[542];
	assign cj_6144[3827] = ci_6144[133];
	assign cj_6144[3828] = ci_6144[684];
	assign cj_6144[3829] = ci_6144[2195];
	assign cj_6144[3830] = ci_6144[4666];
	assign cj_6144[3831] = ci_6144[1953];
	assign cj_6144[3832] = ci_6144[200];
	assign cj_6144[3833] = ci_6144[5551];
	assign cj_6144[3834] = ci_6144[5718];
	assign cj_6144[3835] = ci_6144[701];
	assign cj_6144[3836] = ci_6144[2788];
	assign cj_6144[3837] = ci_6144[5835];
	assign cj_6144[3838] = ci_6144[3698];
	assign cj_6144[3839] = ci_6144[2521];
	assign cj_6144[3840] = ci_6144[2304];
	assign cj_6144[3841] = ci_6144[3047];
	assign cj_6144[3842] = ci_6144[4750];
	assign cj_6144[3843] = ci_6144[1269];
	assign cj_6144[3844] = ci_6144[4892];
	assign cj_6144[3845] = ci_6144[3331];
	assign cj_6144[3846] = ci_6144[2730];
	assign cj_6144[3847] = ci_6144[3089];
	assign cj_6144[3848] = ci_6144[4408];
	assign cj_6144[3849] = ci_6144[543];
	assign cj_6144[3850] = ci_6144[3782];
	assign cj_6144[3851] = ci_6144[1837];
	assign cj_6144[3852] = ci_6144[852];
	assign cj_6144[3853] = ci_6144[827];
	assign cj_6144[3854] = ci_6144[1762];
	assign cj_6144[3855] = ci_6144[3657];
	assign cj_6144[3856] = ci_6144[368];
	assign cj_6144[3857] = ci_6144[4183];
	assign cj_6144[3858] = ci_6144[2814];
	assign cj_6144[3859] = ci_6144[2405];
	assign cj_6144[3860] = ci_6144[2956];
	assign cj_6144[3861] = ci_6144[4467];
	assign cj_6144[3862] = ci_6144[794];
	assign cj_6144[3863] = ci_6144[4225];
	assign cj_6144[3864] = ci_6144[2472];
	assign cj_6144[3865] = ci_6144[1679];
	assign cj_6144[3866] = ci_6144[1846];
	assign cj_6144[3867] = ci_6144[2973];
	assign cj_6144[3868] = ci_6144[5060];
	assign cj_6144[3869] = ci_6144[1963];
	assign cj_6144[3870] = ci_6144[5970];
	assign cj_6144[3871] = ci_6144[4793];
	assign cj_6144[3872] = ci_6144[4576];
	assign cj_6144[3873] = ci_6144[5319];
	assign cj_6144[3874] = ci_6144[878];
	assign cj_6144[3875] = ci_6144[3541];
	assign cj_6144[3876] = ci_6144[1020];
	assign cj_6144[3877] = ci_6144[5603];
	assign cj_6144[3878] = ci_6144[5002];
	assign cj_6144[3879] = ci_6144[5361];
	assign cj_6144[3880] = ci_6144[536];
	assign cj_6144[3881] = ci_6144[2815];
	assign cj_6144[3882] = ci_6144[6054];
	assign cj_6144[3883] = ci_6144[4109];
	assign cj_6144[3884] = ci_6144[3124];
	assign cj_6144[3885] = ci_6144[3099];
	assign cj_6144[3886] = ci_6144[4034];
	assign cj_6144[3887] = ci_6144[5929];
	assign cj_6144[3888] = ci_6144[2640];
	assign cj_6144[3889] = ci_6144[311];
	assign cj_6144[3890] = ci_6144[5086];
	assign cj_6144[3891] = ci_6144[4677];
	assign cj_6144[3892] = ci_6144[5228];
	assign cj_6144[3893] = ci_6144[595];
	assign cj_6144[3894] = ci_6144[3066];
	assign cj_6144[3895] = ci_6144[353];
	assign cj_6144[3896] = ci_6144[4744];
	assign cj_6144[3897] = ci_6144[3951];
	assign cj_6144[3898] = ci_6144[4118];
	assign cj_6144[3899] = ci_6144[5245];
	assign cj_6144[3900] = ci_6144[1188];
	assign cj_6144[3901] = ci_6144[4235];
	assign cj_6144[3902] = ci_6144[2098];
	assign cj_6144[3903] = ci_6144[921];
	assign cj_6144[3904] = ci_6144[704];
	assign cj_6144[3905] = ci_6144[1447];
	assign cj_6144[3906] = ci_6144[3150];
	assign cj_6144[3907] = ci_6144[5813];
	assign cj_6144[3908] = ci_6144[3292];
	assign cj_6144[3909] = ci_6144[1731];
	assign cj_6144[3910] = ci_6144[1130];
	assign cj_6144[3911] = ci_6144[1489];
	assign cj_6144[3912] = ci_6144[2808];
	assign cj_6144[3913] = ci_6144[5087];
	assign cj_6144[3914] = ci_6144[2182];
	assign cj_6144[3915] = ci_6144[237];
	assign cj_6144[3916] = ci_6144[5396];
	assign cj_6144[3917] = ci_6144[5371];
	assign cj_6144[3918] = ci_6144[162];
	assign cj_6144[3919] = ci_6144[2057];
	assign cj_6144[3920] = ci_6144[4912];
	assign cj_6144[3921] = ci_6144[2583];
	assign cj_6144[3922] = ci_6144[1214];
	assign cj_6144[3923] = ci_6144[805];
	assign cj_6144[3924] = ci_6144[1356];
	assign cj_6144[3925] = ci_6144[2867];
	assign cj_6144[3926] = ci_6144[5338];
	assign cj_6144[3927] = ci_6144[2625];
	assign cj_6144[3928] = ci_6144[872];
	assign cj_6144[3929] = ci_6144[79];
	assign cj_6144[3930] = ci_6144[246];
	assign cj_6144[3931] = ci_6144[1373];
	assign cj_6144[3932] = ci_6144[3460];
	assign cj_6144[3933] = ci_6144[363];
	assign cj_6144[3934] = ci_6144[4370];
	assign cj_6144[3935] = ci_6144[3193];
	assign cj_6144[3936] = ci_6144[2976];
	assign cj_6144[3937] = ci_6144[3719];
	assign cj_6144[3938] = ci_6144[5422];
	assign cj_6144[3939] = ci_6144[1941];
	assign cj_6144[3940] = ci_6144[5564];
	assign cj_6144[3941] = ci_6144[4003];
	assign cj_6144[3942] = ci_6144[3402];
	assign cj_6144[3943] = ci_6144[3761];
	assign cj_6144[3944] = ci_6144[5080];
	assign cj_6144[3945] = ci_6144[1215];
	assign cj_6144[3946] = ci_6144[4454];
	assign cj_6144[3947] = ci_6144[2509];
	assign cj_6144[3948] = ci_6144[1524];
	assign cj_6144[3949] = ci_6144[1499];
	assign cj_6144[3950] = ci_6144[2434];
	assign cj_6144[3951] = ci_6144[4329];
	assign cj_6144[3952] = ci_6144[1040];
	assign cj_6144[3953] = ci_6144[4855];
	assign cj_6144[3954] = ci_6144[3486];
	assign cj_6144[3955] = ci_6144[3077];
	assign cj_6144[3956] = ci_6144[3628];
	assign cj_6144[3957] = ci_6144[5139];
	assign cj_6144[3958] = ci_6144[1466];
	assign cj_6144[3959] = ci_6144[4897];
	assign cj_6144[3960] = ci_6144[3144];
	assign cj_6144[3961] = ci_6144[2351];
	assign cj_6144[3962] = ci_6144[2518];
	assign cj_6144[3963] = ci_6144[3645];
	assign cj_6144[3964] = ci_6144[5732];
	assign cj_6144[3965] = ci_6144[2635];
	assign cj_6144[3966] = ci_6144[498];
	assign cj_6144[3967] = ci_6144[5465];
	assign cj_6144[3968] = ci_6144[5248];
	assign cj_6144[3969] = ci_6144[5991];
	assign cj_6144[3970] = ci_6144[1550];
	assign cj_6144[3971] = ci_6144[4213];
	assign cj_6144[3972] = ci_6144[1692];
	assign cj_6144[3973] = ci_6144[131];
	assign cj_6144[3974] = ci_6144[5674];
	assign cj_6144[3975] = ci_6144[6033];
	assign cj_6144[3976] = ci_6144[1208];
	assign cj_6144[3977] = ci_6144[3487];
	assign cj_6144[3978] = ci_6144[582];
	assign cj_6144[3979] = ci_6144[4781];
	assign cj_6144[3980] = ci_6144[3796];
	assign cj_6144[3981] = ci_6144[3771];
	assign cj_6144[3982] = ci_6144[4706];
	assign cj_6144[3983] = ci_6144[457];
	assign cj_6144[3984] = ci_6144[3312];
	assign cj_6144[3985] = ci_6144[983];
	assign cj_6144[3986] = ci_6144[5758];
	assign cj_6144[3987] = ci_6144[5349];
	assign cj_6144[3988] = ci_6144[5900];
	assign cj_6144[3989] = ci_6144[1267];
	assign cj_6144[3990] = ci_6144[3738];
	assign cj_6144[3991] = ci_6144[1025];
	assign cj_6144[3992] = ci_6144[5416];
	assign cj_6144[3993] = ci_6144[4623];
	assign cj_6144[3994] = ci_6144[4790];
	assign cj_6144[3995] = ci_6144[5917];
	assign cj_6144[3996] = ci_6144[1860];
	assign cj_6144[3997] = ci_6144[4907];
	assign cj_6144[3998] = ci_6144[2770];
	assign cj_6144[3999] = ci_6144[1593];
	assign cj_6144[4000] = ci_6144[1376];
	assign cj_6144[4001] = ci_6144[2119];
	assign cj_6144[4002] = ci_6144[3822];
	assign cj_6144[4003] = ci_6144[341];
	assign cj_6144[4004] = ci_6144[3964];
	assign cj_6144[4005] = ci_6144[2403];
	assign cj_6144[4006] = ci_6144[1802];
	assign cj_6144[4007] = ci_6144[2161];
	assign cj_6144[4008] = ci_6144[3480];
	assign cj_6144[4009] = ci_6144[5759];
	assign cj_6144[4010] = ci_6144[2854];
	assign cj_6144[4011] = ci_6144[909];
	assign cj_6144[4012] = ci_6144[6068];
	assign cj_6144[4013] = ci_6144[6043];
	assign cj_6144[4014] = ci_6144[834];
	assign cj_6144[4015] = ci_6144[2729];
	assign cj_6144[4016] = ci_6144[5584];
	assign cj_6144[4017] = ci_6144[3255];
	assign cj_6144[4018] = ci_6144[1886];
	assign cj_6144[4019] = ci_6144[1477];
	assign cj_6144[4020] = ci_6144[2028];
	assign cj_6144[4021] = ci_6144[3539];
	assign cj_6144[4022] = ci_6144[6010];
	assign cj_6144[4023] = ci_6144[3297];
	assign cj_6144[4024] = ci_6144[1544];
	assign cj_6144[4025] = ci_6144[751];
	assign cj_6144[4026] = ci_6144[918];
	assign cj_6144[4027] = ci_6144[2045];
	assign cj_6144[4028] = ci_6144[4132];
	assign cj_6144[4029] = ci_6144[1035];
	assign cj_6144[4030] = ci_6144[5042];
	assign cj_6144[4031] = ci_6144[3865];
	assign cj_6144[4032] = ci_6144[3648];
	assign cj_6144[4033] = ci_6144[4391];
	assign cj_6144[4034] = ci_6144[6094];
	assign cj_6144[4035] = ci_6144[2613];
	assign cj_6144[4036] = ci_6144[92];
	assign cj_6144[4037] = ci_6144[4675];
	assign cj_6144[4038] = ci_6144[4074];
	assign cj_6144[4039] = ci_6144[4433];
	assign cj_6144[4040] = ci_6144[5752];
	assign cj_6144[4041] = ci_6144[1887];
	assign cj_6144[4042] = ci_6144[5126];
	assign cj_6144[4043] = ci_6144[3181];
	assign cj_6144[4044] = ci_6144[2196];
	assign cj_6144[4045] = ci_6144[2171];
	assign cj_6144[4046] = ci_6144[3106];
	assign cj_6144[4047] = ci_6144[5001];
	assign cj_6144[4048] = ci_6144[1712];
	assign cj_6144[4049] = ci_6144[5527];
	assign cj_6144[4050] = ci_6144[4158];
	assign cj_6144[4051] = ci_6144[3749];
	assign cj_6144[4052] = ci_6144[4300];
	assign cj_6144[4053] = ci_6144[5811];
	assign cj_6144[4054] = ci_6144[2138];
	assign cj_6144[4055] = ci_6144[5569];
	assign cj_6144[4056] = ci_6144[3816];
	assign cj_6144[4057] = ci_6144[3023];
	assign cj_6144[4058] = ci_6144[3190];
	assign cj_6144[4059] = ci_6144[4317];
	assign cj_6144[4060] = ci_6144[260];
	assign cj_6144[4061] = ci_6144[3307];
	assign cj_6144[4062] = ci_6144[1170];
	assign cj_6144[4063] = ci_6144[6137];
	assign cj_6144[4064] = ci_6144[5920];
	assign cj_6144[4065] = ci_6144[519];
	assign cj_6144[4066] = ci_6144[2222];
	assign cj_6144[4067] = ci_6144[4885];
	assign cj_6144[4068] = ci_6144[2364];
	assign cj_6144[4069] = ci_6144[803];
	assign cj_6144[4070] = ci_6144[202];
	assign cj_6144[4071] = ci_6144[561];
	assign cj_6144[4072] = ci_6144[1880];
	assign cj_6144[4073] = ci_6144[4159];
	assign cj_6144[4074] = ci_6144[1254];
	assign cj_6144[4075] = ci_6144[5453];
	assign cj_6144[4076] = ci_6144[4468];
	assign cj_6144[4077] = ci_6144[4443];
	assign cj_6144[4078] = ci_6144[5378];
	assign cj_6144[4079] = ci_6144[1129];
	assign cj_6144[4080] = ci_6144[3984];
	assign cj_6144[4081] = ci_6144[1655];
	assign cj_6144[4082] = ci_6144[286];
	assign cj_6144[4083] = ci_6144[6021];
	assign cj_6144[4084] = ci_6144[428];
	assign cj_6144[4085] = ci_6144[1939];
	assign cj_6144[4086] = ci_6144[4410];
	assign cj_6144[4087] = ci_6144[1697];
	assign cj_6144[4088] = ci_6144[6088];
	assign cj_6144[4089] = ci_6144[5295];
	assign cj_6144[4090] = ci_6144[5462];
	assign cj_6144[4091] = ci_6144[445];
	assign cj_6144[4092] = ci_6144[2532];
	assign cj_6144[4093] = ci_6144[5579];
	assign cj_6144[4094] = ci_6144[3442];
	assign cj_6144[4095] = ci_6144[2265];
	assign cj_6144[4096] = ci_6144[2048];
	assign cj_6144[4097] = ci_6144[2791];
	assign cj_6144[4098] = ci_6144[4494];
	assign cj_6144[4099] = ci_6144[1013];
	assign cj_6144[4100] = ci_6144[4636];
	assign cj_6144[4101] = ci_6144[3075];
	assign cj_6144[4102] = ci_6144[2474];
	assign cj_6144[4103] = ci_6144[2833];
	assign cj_6144[4104] = ci_6144[4152];
	assign cj_6144[4105] = ci_6144[287];
	assign cj_6144[4106] = ci_6144[3526];
	assign cj_6144[4107] = ci_6144[1581];
	assign cj_6144[4108] = ci_6144[596];
	assign cj_6144[4109] = ci_6144[571];
	assign cj_6144[4110] = ci_6144[1506];
	assign cj_6144[4111] = ci_6144[3401];
	assign cj_6144[4112] = ci_6144[112];
	assign cj_6144[4113] = ci_6144[3927];
	assign cj_6144[4114] = ci_6144[2558];
	assign cj_6144[4115] = ci_6144[2149];
	assign cj_6144[4116] = ci_6144[2700];
	assign cj_6144[4117] = ci_6144[4211];
	assign cj_6144[4118] = ci_6144[538];
	assign cj_6144[4119] = ci_6144[3969];
	assign cj_6144[4120] = ci_6144[2216];
	assign cj_6144[4121] = ci_6144[1423];
	assign cj_6144[4122] = ci_6144[1590];
	assign cj_6144[4123] = ci_6144[2717];
	assign cj_6144[4124] = ci_6144[4804];
	assign cj_6144[4125] = ci_6144[1707];
	assign cj_6144[4126] = ci_6144[5714];
	assign cj_6144[4127] = ci_6144[4537];
	assign cj_6144[4128] = ci_6144[4320];
	assign cj_6144[4129] = ci_6144[5063];
	assign cj_6144[4130] = ci_6144[622];
	assign cj_6144[4131] = ci_6144[3285];
	assign cj_6144[4132] = ci_6144[764];
	assign cj_6144[4133] = ci_6144[5347];
	assign cj_6144[4134] = ci_6144[4746];
	assign cj_6144[4135] = ci_6144[5105];
	assign cj_6144[4136] = ci_6144[280];
	assign cj_6144[4137] = ci_6144[2559];
	assign cj_6144[4138] = ci_6144[5798];
	assign cj_6144[4139] = ci_6144[3853];
	assign cj_6144[4140] = ci_6144[2868];
	assign cj_6144[4141] = ci_6144[2843];
	assign cj_6144[4142] = ci_6144[3778];
	assign cj_6144[4143] = ci_6144[5673];
	assign cj_6144[4144] = ci_6144[2384];
	assign cj_6144[4145] = ci_6144[55];
	assign cj_6144[4146] = ci_6144[4830];
	assign cj_6144[4147] = ci_6144[4421];
	assign cj_6144[4148] = ci_6144[4972];
	assign cj_6144[4149] = ci_6144[339];
	assign cj_6144[4150] = ci_6144[2810];
	assign cj_6144[4151] = ci_6144[97];
	assign cj_6144[4152] = ci_6144[4488];
	assign cj_6144[4153] = ci_6144[3695];
	assign cj_6144[4154] = ci_6144[3862];
	assign cj_6144[4155] = ci_6144[4989];
	assign cj_6144[4156] = ci_6144[932];
	assign cj_6144[4157] = ci_6144[3979];
	assign cj_6144[4158] = ci_6144[1842];
	assign cj_6144[4159] = ci_6144[665];
	assign cj_6144[4160] = ci_6144[448];
	assign cj_6144[4161] = ci_6144[1191];
	assign cj_6144[4162] = ci_6144[2894];
	assign cj_6144[4163] = ci_6144[5557];
	assign cj_6144[4164] = ci_6144[3036];
	assign cj_6144[4165] = ci_6144[1475];
	assign cj_6144[4166] = ci_6144[874];
	assign cj_6144[4167] = ci_6144[1233];
	assign cj_6144[4168] = ci_6144[2552];
	assign cj_6144[4169] = ci_6144[4831];
	assign cj_6144[4170] = ci_6144[1926];
	assign cj_6144[4171] = ci_6144[6125];
	assign cj_6144[4172] = ci_6144[5140];
	assign cj_6144[4173] = ci_6144[5115];
	assign cj_6144[4174] = ci_6144[6050];
	assign cj_6144[4175] = ci_6144[1801];
	assign cj_6144[4176] = ci_6144[4656];
	assign cj_6144[4177] = ci_6144[2327];
	assign cj_6144[4178] = ci_6144[958];
	assign cj_6144[4179] = ci_6144[549];
	assign cj_6144[4180] = ci_6144[1100];
	assign cj_6144[4181] = ci_6144[2611];
	assign cj_6144[4182] = ci_6144[5082];
	assign cj_6144[4183] = ci_6144[2369];
	assign cj_6144[4184] = ci_6144[616];
	assign cj_6144[4185] = ci_6144[5967];
	assign cj_6144[4186] = ci_6144[6134];
	assign cj_6144[4187] = ci_6144[1117];
	assign cj_6144[4188] = ci_6144[3204];
	assign cj_6144[4189] = ci_6144[107];
	assign cj_6144[4190] = ci_6144[4114];
	assign cj_6144[4191] = ci_6144[2937];
	assign cj_6144[4192] = ci_6144[2720];
	assign cj_6144[4193] = ci_6144[3463];
	assign cj_6144[4194] = ci_6144[5166];
	assign cj_6144[4195] = ci_6144[1685];
	assign cj_6144[4196] = ci_6144[5308];
	assign cj_6144[4197] = ci_6144[3747];
	assign cj_6144[4198] = ci_6144[3146];
	assign cj_6144[4199] = ci_6144[3505];
	assign cj_6144[4200] = ci_6144[4824];
	assign cj_6144[4201] = ci_6144[959];
	assign cj_6144[4202] = ci_6144[4198];
	assign cj_6144[4203] = ci_6144[2253];
	assign cj_6144[4204] = ci_6144[1268];
	assign cj_6144[4205] = ci_6144[1243];
	assign cj_6144[4206] = ci_6144[2178];
	assign cj_6144[4207] = ci_6144[4073];
	assign cj_6144[4208] = ci_6144[784];
	assign cj_6144[4209] = ci_6144[4599];
	assign cj_6144[4210] = ci_6144[3230];
	assign cj_6144[4211] = ci_6144[2821];
	assign cj_6144[4212] = ci_6144[3372];
	assign cj_6144[4213] = ci_6144[4883];
	assign cj_6144[4214] = ci_6144[1210];
	assign cj_6144[4215] = ci_6144[4641];
	assign cj_6144[4216] = ci_6144[2888];
	assign cj_6144[4217] = ci_6144[2095];
	assign cj_6144[4218] = ci_6144[2262];
	assign cj_6144[4219] = ci_6144[3389];
	assign cj_6144[4220] = ci_6144[5476];
	assign cj_6144[4221] = ci_6144[2379];
	assign cj_6144[4222] = ci_6144[242];
	assign cj_6144[4223] = ci_6144[5209];
	assign cj_6144[4224] = ci_6144[4992];
	assign cj_6144[4225] = ci_6144[5735];
	assign cj_6144[4226] = ci_6144[1294];
	assign cj_6144[4227] = ci_6144[3957];
	assign cj_6144[4228] = ci_6144[1436];
	assign cj_6144[4229] = ci_6144[6019];
	assign cj_6144[4230] = ci_6144[5418];
	assign cj_6144[4231] = ci_6144[5777];
	assign cj_6144[4232] = ci_6144[952];
	assign cj_6144[4233] = ci_6144[3231];
	assign cj_6144[4234] = ci_6144[326];
	assign cj_6144[4235] = ci_6144[4525];
	assign cj_6144[4236] = ci_6144[3540];
	assign cj_6144[4237] = ci_6144[3515];
	assign cj_6144[4238] = ci_6144[4450];
	assign cj_6144[4239] = ci_6144[201];
	assign cj_6144[4240] = ci_6144[3056];
	assign cj_6144[4241] = ci_6144[727];
	assign cj_6144[4242] = ci_6144[5502];
	assign cj_6144[4243] = ci_6144[5093];
	assign cj_6144[4244] = ci_6144[5644];
	assign cj_6144[4245] = ci_6144[1011];
	assign cj_6144[4246] = ci_6144[3482];
	assign cj_6144[4247] = ci_6144[769];
	assign cj_6144[4248] = ci_6144[5160];
	assign cj_6144[4249] = ci_6144[4367];
	assign cj_6144[4250] = ci_6144[4534];
	assign cj_6144[4251] = ci_6144[5661];
	assign cj_6144[4252] = ci_6144[1604];
	assign cj_6144[4253] = ci_6144[4651];
	assign cj_6144[4254] = ci_6144[2514];
	assign cj_6144[4255] = ci_6144[1337];
	assign cj_6144[4256] = ci_6144[1120];
	assign cj_6144[4257] = ci_6144[1863];
	assign cj_6144[4258] = ci_6144[3566];
	assign cj_6144[4259] = ci_6144[85];
	assign cj_6144[4260] = ci_6144[3708];
	assign cj_6144[4261] = ci_6144[2147];
	assign cj_6144[4262] = ci_6144[1546];
	assign cj_6144[4263] = ci_6144[1905];
	assign cj_6144[4264] = ci_6144[3224];
	assign cj_6144[4265] = ci_6144[5503];
	assign cj_6144[4266] = ci_6144[2598];
	assign cj_6144[4267] = ci_6144[653];
	assign cj_6144[4268] = ci_6144[5812];
	assign cj_6144[4269] = ci_6144[5787];
	assign cj_6144[4270] = ci_6144[578];
	assign cj_6144[4271] = ci_6144[2473];
	assign cj_6144[4272] = ci_6144[5328];
	assign cj_6144[4273] = ci_6144[2999];
	assign cj_6144[4274] = ci_6144[1630];
	assign cj_6144[4275] = ci_6144[1221];
	assign cj_6144[4276] = ci_6144[1772];
	assign cj_6144[4277] = ci_6144[3283];
	assign cj_6144[4278] = ci_6144[5754];
	assign cj_6144[4279] = ci_6144[3041];
	assign cj_6144[4280] = ci_6144[1288];
	assign cj_6144[4281] = ci_6144[495];
	assign cj_6144[4282] = ci_6144[662];
	assign cj_6144[4283] = ci_6144[1789];
	assign cj_6144[4284] = ci_6144[3876];
	assign cj_6144[4285] = ci_6144[779];
	assign cj_6144[4286] = ci_6144[4786];
	assign cj_6144[4287] = ci_6144[3609];
	assign cj_6144[4288] = ci_6144[3392];
	assign cj_6144[4289] = ci_6144[4135];
	assign cj_6144[4290] = ci_6144[5838];
	assign cj_6144[4291] = ci_6144[2357];
	assign cj_6144[4292] = ci_6144[5980];
	assign cj_6144[4293] = ci_6144[4419];
	assign cj_6144[4294] = ci_6144[3818];
	assign cj_6144[4295] = ci_6144[4177];
	assign cj_6144[4296] = ci_6144[5496];
	assign cj_6144[4297] = ci_6144[1631];
	assign cj_6144[4298] = ci_6144[4870];
	assign cj_6144[4299] = ci_6144[2925];
	assign cj_6144[4300] = ci_6144[1940];
	assign cj_6144[4301] = ci_6144[1915];
	assign cj_6144[4302] = ci_6144[2850];
	assign cj_6144[4303] = ci_6144[4745];
	assign cj_6144[4304] = ci_6144[1456];
	assign cj_6144[4305] = ci_6144[5271];
	assign cj_6144[4306] = ci_6144[3902];
	assign cj_6144[4307] = ci_6144[3493];
	assign cj_6144[4308] = ci_6144[4044];
	assign cj_6144[4309] = ci_6144[5555];
	assign cj_6144[4310] = ci_6144[1882];
	assign cj_6144[4311] = ci_6144[5313];
	assign cj_6144[4312] = ci_6144[3560];
	assign cj_6144[4313] = ci_6144[2767];
	assign cj_6144[4314] = ci_6144[2934];
	assign cj_6144[4315] = ci_6144[4061];
	assign cj_6144[4316] = ci_6144[4];
	assign cj_6144[4317] = ci_6144[3051];
	assign cj_6144[4318] = ci_6144[914];
	assign cj_6144[4319] = ci_6144[5881];
	assign cj_6144[4320] = ci_6144[5664];
	assign cj_6144[4321] = ci_6144[263];
	assign cj_6144[4322] = ci_6144[1966];
	assign cj_6144[4323] = ci_6144[4629];
	assign cj_6144[4324] = ci_6144[2108];
	assign cj_6144[4325] = ci_6144[547];
	assign cj_6144[4326] = ci_6144[6090];
	assign cj_6144[4327] = ci_6144[305];
	assign cj_6144[4328] = ci_6144[1624];
	assign cj_6144[4329] = ci_6144[3903];
	assign cj_6144[4330] = ci_6144[998];
	assign cj_6144[4331] = ci_6144[5197];
	assign cj_6144[4332] = ci_6144[4212];
	assign cj_6144[4333] = ci_6144[4187];
	assign cj_6144[4334] = ci_6144[5122];
	assign cj_6144[4335] = ci_6144[873];
	assign cj_6144[4336] = ci_6144[3728];
	assign cj_6144[4337] = ci_6144[1399];
	assign cj_6144[4338] = ci_6144[30];
	assign cj_6144[4339] = ci_6144[5765];
	assign cj_6144[4340] = ci_6144[172];
	assign cj_6144[4341] = ci_6144[1683];
	assign cj_6144[4342] = ci_6144[4154];
	assign cj_6144[4343] = ci_6144[1441];
	assign cj_6144[4344] = ci_6144[5832];
	assign cj_6144[4345] = ci_6144[5039];
	assign cj_6144[4346] = ci_6144[5206];
	assign cj_6144[4347] = ci_6144[189];
	assign cj_6144[4348] = ci_6144[2276];
	assign cj_6144[4349] = ci_6144[5323];
	assign cj_6144[4350] = ci_6144[3186];
	assign cj_6144[4351] = ci_6144[2009];
	assign cj_6144[4352] = ci_6144[1792];
	assign cj_6144[4353] = ci_6144[2535];
	assign cj_6144[4354] = ci_6144[4238];
	assign cj_6144[4355] = ci_6144[757];
	assign cj_6144[4356] = ci_6144[4380];
	assign cj_6144[4357] = ci_6144[2819];
	assign cj_6144[4358] = ci_6144[2218];
	assign cj_6144[4359] = ci_6144[2577];
	assign cj_6144[4360] = ci_6144[3896];
	assign cj_6144[4361] = ci_6144[31];
	assign cj_6144[4362] = ci_6144[3270];
	assign cj_6144[4363] = ci_6144[1325];
	assign cj_6144[4364] = ci_6144[340];
	assign cj_6144[4365] = ci_6144[315];
	assign cj_6144[4366] = ci_6144[1250];
	assign cj_6144[4367] = ci_6144[3145];
	assign cj_6144[4368] = ci_6144[6000];
	assign cj_6144[4369] = ci_6144[3671];
	assign cj_6144[4370] = ci_6144[2302];
	assign cj_6144[4371] = ci_6144[1893];
	assign cj_6144[4372] = ci_6144[2444];
	assign cj_6144[4373] = ci_6144[3955];
	assign cj_6144[4374] = ci_6144[282];
	assign cj_6144[4375] = ci_6144[3713];
	assign cj_6144[4376] = ci_6144[1960];
	assign cj_6144[4377] = ci_6144[1167];
	assign cj_6144[4378] = ci_6144[1334];
	assign cj_6144[4379] = ci_6144[2461];
	assign cj_6144[4380] = ci_6144[4548];
	assign cj_6144[4381] = ci_6144[1451];
	assign cj_6144[4382] = ci_6144[5458];
	assign cj_6144[4383] = ci_6144[4281];
	assign cj_6144[4384] = ci_6144[4064];
	assign cj_6144[4385] = ci_6144[4807];
	assign cj_6144[4386] = ci_6144[366];
	assign cj_6144[4387] = ci_6144[3029];
	assign cj_6144[4388] = ci_6144[508];
	assign cj_6144[4389] = ci_6144[5091];
	assign cj_6144[4390] = ci_6144[4490];
	assign cj_6144[4391] = ci_6144[4849];
	assign cj_6144[4392] = ci_6144[24];
	assign cj_6144[4393] = ci_6144[2303];
	assign cj_6144[4394] = ci_6144[5542];
	assign cj_6144[4395] = ci_6144[3597];
	assign cj_6144[4396] = ci_6144[2612];
	assign cj_6144[4397] = ci_6144[2587];
	assign cj_6144[4398] = ci_6144[3522];
	assign cj_6144[4399] = ci_6144[5417];
	assign cj_6144[4400] = ci_6144[2128];
	assign cj_6144[4401] = ci_6144[5943];
	assign cj_6144[4402] = ci_6144[4574];
	assign cj_6144[4403] = ci_6144[4165];
	assign cj_6144[4404] = ci_6144[4716];
	assign cj_6144[4405] = ci_6144[83];
	assign cj_6144[4406] = ci_6144[2554];
	assign cj_6144[4407] = ci_6144[5985];
	assign cj_6144[4408] = ci_6144[4232];
	assign cj_6144[4409] = ci_6144[3439];
	assign cj_6144[4410] = ci_6144[3606];
	assign cj_6144[4411] = ci_6144[4733];
	assign cj_6144[4412] = ci_6144[676];
	assign cj_6144[4413] = ci_6144[3723];
	assign cj_6144[4414] = ci_6144[1586];
	assign cj_6144[4415] = ci_6144[409];
	assign cj_6144[4416] = ci_6144[192];
	assign cj_6144[4417] = ci_6144[935];
	assign cj_6144[4418] = ci_6144[2638];
	assign cj_6144[4419] = ci_6144[5301];
	assign cj_6144[4420] = ci_6144[2780];
	assign cj_6144[4421] = ci_6144[1219];
	assign cj_6144[4422] = ci_6144[618];
	assign cj_6144[4423] = ci_6144[977];
	assign cj_6144[4424] = ci_6144[2296];
	assign cj_6144[4425] = ci_6144[4575];
	assign cj_6144[4426] = ci_6144[1670];
	assign cj_6144[4427] = ci_6144[5869];
	assign cj_6144[4428] = ci_6144[4884];
	assign cj_6144[4429] = ci_6144[4859];
	assign cj_6144[4430] = ci_6144[5794];
	assign cj_6144[4431] = ci_6144[1545];
	assign cj_6144[4432] = ci_6144[4400];
	assign cj_6144[4433] = ci_6144[2071];
	assign cj_6144[4434] = ci_6144[702];
	assign cj_6144[4435] = ci_6144[293];
	assign cj_6144[4436] = ci_6144[844];
	assign cj_6144[4437] = ci_6144[2355];
	assign cj_6144[4438] = ci_6144[4826];
	assign cj_6144[4439] = ci_6144[2113];
	assign cj_6144[4440] = ci_6144[360];
	assign cj_6144[4441] = ci_6144[5711];
	assign cj_6144[4442] = ci_6144[5878];
	assign cj_6144[4443] = ci_6144[861];
	assign cj_6144[4444] = ci_6144[2948];
	assign cj_6144[4445] = ci_6144[5995];
	assign cj_6144[4446] = ci_6144[3858];
	assign cj_6144[4447] = ci_6144[2681];
	assign cj_6144[4448] = ci_6144[2464];
	assign cj_6144[4449] = ci_6144[3207];
	assign cj_6144[4450] = ci_6144[4910];
	assign cj_6144[4451] = ci_6144[1429];
	assign cj_6144[4452] = ci_6144[5052];
	assign cj_6144[4453] = ci_6144[3491];
	assign cj_6144[4454] = ci_6144[2890];
	assign cj_6144[4455] = ci_6144[3249];
	assign cj_6144[4456] = ci_6144[4568];
	assign cj_6144[4457] = ci_6144[703];
	assign cj_6144[4458] = ci_6144[3942];
	assign cj_6144[4459] = ci_6144[1997];
	assign cj_6144[4460] = ci_6144[1012];
	assign cj_6144[4461] = ci_6144[987];
	assign cj_6144[4462] = ci_6144[1922];
	assign cj_6144[4463] = ci_6144[3817];
	assign cj_6144[4464] = ci_6144[528];
	assign cj_6144[4465] = ci_6144[4343];
	assign cj_6144[4466] = ci_6144[2974];
	assign cj_6144[4467] = ci_6144[2565];
	assign cj_6144[4468] = ci_6144[3116];
	assign cj_6144[4469] = ci_6144[4627];
	assign cj_6144[4470] = ci_6144[954];
	assign cj_6144[4471] = ci_6144[4385];
	assign cj_6144[4472] = ci_6144[2632];
	assign cj_6144[4473] = ci_6144[1839];
	assign cj_6144[4474] = ci_6144[2006];
	assign cj_6144[4475] = ci_6144[3133];
	assign cj_6144[4476] = ci_6144[5220];
	assign cj_6144[4477] = ci_6144[2123];
	assign cj_6144[4478] = ci_6144[6130];
	assign cj_6144[4479] = ci_6144[4953];
	assign cj_6144[4480] = ci_6144[4736];
	assign cj_6144[4481] = ci_6144[5479];
	assign cj_6144[4482] = ci_6144[1038];
	assign cj_6144[4483] = ci_6144[3701];
	assign cj_6144[4484] = ci_6144[1180];
	assign cj_6144[4485] = ci_6144[5763];
	assign cj_6144[4486] = ci_6144[5162];
	assign cj_6144[4487] = ci_6144[5521];
	assign cj_6144[4488] = ci_6144[696];
	assign cj_6144[4489] = ci_6144[2975];
	assign cj_6144[4490] = ci_6144[70];
	assign cj_6144[4491] = ci_6144[4269];
	assign cj_6144[4492] = ci_6144[3284];
	assign cj_6144[4493] = ci_6144[3259];
	assign cj_6144[4494] = ci_6144[4194];
	assign cj_6144[4495] = ci_6144[6089];
	assign cj_6144[4496] = ci_6144[2800];
	assign cj_6144[4497] = ci_6144[471];
	assign cj_6144[4498] = ci_6144[5246];
	assign cj_6144[4499] = ci_6144[4837];
	assign cj_6144[4500] = ci_6144[5388];
	assign cj_6144[4501] = ci_6144[755];
	assign cj_6144[4502] = ci_6144[3226];
	assign cj_6144[4503] = ci_6144[513];
	assign cj_6144[4504] = ci_6144[4904];
	assign cj_6144[4505] = ci_6144[4111];
	assign cj_6144[4506] = ci_6144[4278];
	assign cj_6144[4507] = ci_6144[5405];
	assign cj_6144[4508] = ci_6144[1348];
	assign cj_6144[4509] = ci_6144[4395];
	assign cj_6144[4510] = ci_6144[2258];
	assign cj_6144[4511] = ci_6144[1081];
	assign cj_6144[4512] = ci_6144[864];
	assign cj_6144[4513] = ci_6144[1607];
	assign cj_6144[4514] = ci_6144[3310];
	assign cj_6144[4515] = ci_6144[5973];
	assign cj_6144[4516] = ci_6144[3452];
	assign cj_6144[4517] = ci_6144[1891];
	assign cj_6144[4518] = ci_6144[1290];
	assign cj_6144[4519] = ci_6144[1649];
	assign cj_6144[4520] = ci_6144[2968];
	assign cj_6144[4521] = ci_6144[5247];
	assign cj_6144[4522] = ci_6144[2342];
	assign cj_6144[4523] = ci_6144[397];
	assign cj_6144[4524] = ci_6144[5556];
	assign cj_6144[4525] = ci_6144[5531];
	assign cj_6144[4526] = ci_6144[322];
	assign cj_6144[4527] = ci_6144[2217];
	assign cj_6144[4528] = ci_6144[5072];
	assign cj_6144[4529] = ci_6144[2743];
	assign cj_6144[4530] = ci_6144[1374];
	assign cj_6144[4531] = ci_6144[965];
	assign cj_6144[4532] = ci_6144[1516];
	assign cj_6144[4533] = ci_6144[3027];
	assign cj_6144[4534] = ci_6144[5498];
	assign cj_6144[4535] = ci_6144[2785];
	assign cj_6144[4536] = ci_6144[1032];
	assign cj_6144[4537] = ci_6144[239];
	assign cj_6144[4538] = ci_6144[406];
	assign cj_6144[4539] = ci_6144[1533];
	assign cj_6144[4540] = ci_6144[3620];
	assign cj_6144[4541] = ci_6144[523];
	assign cj_6144[4542] = ci_6144[4530];
	assign cj_6144[4543] = ci_6144[3353];
	assign cj_6144[4544] = ci_6144[3136];
	assign cj_6144[4545] = ci_6144[3879];
	assign cj_6144[4546] = ci_6144[5582];
	assign cj_6144[4547] = ci_6144[2101];
	assign cj_6144[4548] = ci_6144[5724];
	assign cj_6144[4549] = ci_6144[4163];
	assign cj_6144[4550] = ci_6144[3562];
	assign cj_6144[4551] = ci_6144[3921];
	assign cj_6144[4552] = ci_6144[5240];
	assign cj_6144[4553] = ci_6144[1375];
	assign cj_6144[4554] = ci_6144[4614];
	assign cj_6144[4555] = ci_6144[2669];
	assign cj_6144[4556] = ci_6144[1684];
	assign cj_6144[4557] = ci_6144[1659];
	assign cj_6144[4558] = ci_6144[2594];
	assign cj_6144[4559] = ci_6144[4489];
	assign cj_6144[4560] = ci_6144[1200];
	assign cj_6144[4561] = ci_6144[5015];
	assign cj_6144[4562] = ci_6144[3646];
	assign cj_6144[4563] = ci_6144[3237];
	assign cj_6144[4564] = ci_6144[3788];
	assign cj_6144[4565] = ci_6144[5299];
	assign cj_6144[4566] = ci_6144[1626];
	assign cj_6144[4567] = ci_6144[5057];
	assign cj_6144[4568] = ci_6144[3304];
	assign cj_6144[4569] = ci_6144[2511];
	assign cj_6144[4570] = ci_6144[2678];
	assign cj_6144[4571] = ci_6144[3805];
	assign cj_6144[4572] = ci_6144[5892];
	assign cj_6144[4573] = ci_6144[2795];
	assign cj_6144[4574] = ci_6144[658];
	assign cj_6144[4575] = ci_6144[5625];
	assign cj_6144[4576] = ci_6144[5408];
	assign cj_6144[4577] = ci_6144[7];
	assign cj_6144[4578] = ci_6144[1710];
	assign cj_6144[4579] = ci_6144[4373];
	assign cj_6144[4580] = ci_6144[1852];
	assign cj_6144[4581] = ci_6144[291];
	assign cj_6144[4582] = ci_6144[5834];
	assign cj_6144[4583] = ci_6144[49];
	assign cj_6144[4584] = ci_6144[1368];
	assign cj_6144[4585] = ci_6144[3647];
	assign cj_6144[4586] = ci_6144[742];
	assign cj_6144[4587] = ci_6144[4941];
	assign cj_6144[4588] = ci_6144[3956];
	assign cj_6144[4589] = ci_6144[3931];
	assign cj_6144[4590] = ci_6144[4866];
	assign cj_6144[4591] = ci_6144[617];
	assign cj_6144[4592] = ci_6144[3472];
	assign cj_6144[4593] = ci_6144[1143];
	assign cj_6144[4594] = ci_6144[5918];
	assign cj_6144[4595] = ci_6144[5509];
	assign cj_6144[4596] = ci_6144[6060];
	assign cj_6144[4597] = ci_6144[1427];
	assign cj_6144[4598] = ci_6144[3898];
	assign cj_6144[4599] = ci_6144[1185];
	assign cj_6144[4600] = ci_6144[5576];
	assign cj_6144[4601] = ci_6144[4783];
	assign cj_6144[4602] = ci_6144[4950];
	assign cj_6144[4603] = ci_6144[6077];
	assign cj_6144[4604] = ci_6144[2020];
	assign cj_6144[4605] = ci_6144[5067];
	assign cj_6144[4606] = ci_6144[2930];
	assign cj_6144[4607] = ci_6144[1753];
	assign cj_6144[4608] = ci_6144[1536];
	assign cj_6144[4609] = ci_6144[2279];
	assign cj_6144[4610] = ci_6144[3982];
	assign cj_6144[4611] = ci_6144[501];
	assign cj_6144[4612] = ci_6144[4124];
	assign cj_6144[4613] = ci_6144[2563];
	assign cj_6144[4614] = ci_6144[1962];
	assign cj_6144[4615] = ci_6144[2321];
	assign cj_6144[4616] = ci_6144[3640];
	assign cj_6144[4617] = ci_6144[5919];
	assign cj_6144[4618] = ci_6144[3014];
	assign cj_6144[4619] = ci_6144[1069];
	assign cj_6144[4620] = ci_6144[84];
	assign cj_6144[4621] = ci_6144[59];
	assign cj_6144[4622] = ci_6144[994];
	assign cj_6144[4623] = ci_6144[2889];
	assign cj_6144[4624] = ci_6144[5744];
	assign cj_6144[4625] = ci_6144[3415];
	assign cj_6144[4626] = ci_6144[2046];
	assign cj_6144[4627] = ci_6144[1637];
	assign cj_6144[4628] = ci_6144[2188];
	assign cj_6144[4629] = ci_6144[3699];
	assign cj_6144[4630] = ci_6144[26];
	assign cj_6144[4631] = ci_6144[3457];
	assign cj_6144[4632] = ci_6144[1704];
	assign cj_6144[4633] = ci_6144[911];
	assign cj_6144[4634] = ci_6144[1078];
	assign cj_6144[4635] = ci_6144[2205];
	assign cj_6144[4636] = ci_6144[4292];
	assign cj_6144[4637] = ci_6144[1195];
	assign cj_6144[4638] = ci_6144[5202];
	assign cj_6144[4639] = ci_6144[4025];
	assign cj_6144[4640] = ci_6144[3808];
	assign cj_6144[4641] = ci_6144[4551];
	assign cj_6144[4642] = ci_6144[110];
	assign cj_6144[4643] = ci_6144[2773];
	assign cj_6144[4644] = ci_6144[252];
	assign cj_6144[4645] = ci_6144[4835];
	assign cj_6144[4646] = ci_6144[4234];
	assign cj_6144[4647] = ci_6144[4593];
	assign cj_6144[4648] = ci_6144[5912];
	assign cj_6144[4649] = ci_6144[2047];
	assign cj_6144[4650] = ci_6144[5286];
	assign cj_6144[4651] = ci_6144[3341];
	assign cj_6144[4652] = ci_6144[2356];
	assign cj_6144[4653] = ci_6144[2331];
	assign cj_6144[4654] = ci_6144[3266];
	assign cj_6144[4655] = ci_6144[5161];
	assign cj_6144[4656] = ci_6144[1872];
	assign cj_6144[4657] = ci_6144[5687];
	assign cj_6144[4658] = ci_6144[4318];
	assign cj_6144[4659] = ci_6144[3909];
	assign cj_6144[4660] = ci_6144[4460];
	assign cj_6144[4661] = ci_6144[5971];
	assign cj_6144[4662] = ci_6144[2298];
	assign cj_6144[4663] = ci_6144[5729];
	assign cj_6144[4664] = ci_6144[3976];
	assign cj_6144[4665] = ci_6144[3183];
	assign cj_6144[4666] = ci_6144[3350];
	assign cj_6144[4667] = ci_6144[4477];
	assign cj_6144[4668] = ci_6144[420];
	assign cj_6144[4669] = ci_6144[3467];
	assign cj_6144[4670] = ci_6144[1330];
	assign cj_6144[4671] = ci_6144[153];
	assign cj_6144[4672] = ci_6144[6080];
	assign cj_6144[4673] = ci_6144[679];
	assign cj_6144[4674] = ci_6144[2382];
	assign cj_6144[4675] = ci_6144[5045];
	assign cj_6144[4676] = ci_6144[2524];
	assign cj_6144[4677] = ci_6144[963];
	assign cj_6144[4678] = ci_6144[362];
	assign cj_6144[4679] = ci_6144[721];
	assign cj_6144[4680] = ci_6144[2040];
	assign cj_6144[4681] = ci_6144[4319];
	assign cj_6144[4682] = ci_6144[1414];
	assign cj_6144[4683] = ci_6144[5613];
	assign cj_6144[4684] = ci_6144[4628];
	assign cj_6144[4685] = ci_6144[4603];
	assign cj_6144[4686] = ci_6144[5538];
	assign cj_6144[4687] = ci_6144[1289];
	assign cj_6144[4688] = ci_6144[4144];
	assign cj_6144[4689] = ci_6144[1815];
	assign cj_6144[4690] = ci_6144[446];
	assign cj_6144[4691] = ci_6144[37];
	assign cj_6144[4692] = ci_6144[588];
	assign cj_6144[4693] = ci_6144[2099];
	assign cj_6144[4694] = ci_6144[4570];
	assign cj_6144[4695] = ci_6144[1857];
	assign cj_6144[4696] = ci_6144[104];
	assign cj_6144[4697] = ci_6144[5455];
	assign cj_6144[4698] = ci_6144[5622];
	assign cj_6144[4699] = ci_6144[605];
	assign cj_6144[4700] = ci_6144[2692];
	assign cj_6144[4701] = ci_6144[5739];
	assign cj_6144[4702] = ci_6144[3602];
	assign cj_6144[4703] = ci_6144[2425];
	assign cj_6144[4704] = ci_6144[2208];
	assign cj_6144[4705] = ci_6144[2951];
	assign cj_6144[4706] = ci_6144[4654];
	assign cj_6144[4707] = ci_6144[1173];
	assign cj_6144[4708] = ci_6144[4796];
	assign cj_6144[4709] = ci_6144[3235];
	assign cj_6144[4710] = ci_6144[2634];
	assign cj_6144[4711] = ci_6144[2993];
	assign cj_6144[4712] = ci_6144[4312];
	assign cj_6144[4713] = ci_6144[447];
	assign cj_6144[4714] = ci_6144[3686];
	assign cj_6144[4715] = ci_6144[1741];
	assign cj_6144[4716] = ci_6144[756];
	assign cj_6144[4717] = ci_6144[731];
	assign cj_6144[4718] = ci_6144[1666];
	assign cj_6144[4719] = ci_6144[3561];
	assign cj_6144[4720] = ci_6144[272];
	assign cj_6144[4721] = ci_6144[4087];
	assign cj_6144[4722] = ci_6144[2718];
	assign cj_6144[4723] = ci_6144[2309];
	assign cj_6144[4724] = ci_6144[2860];
	assign cj_6144[4725] = ci_6144[4371];
	assign cj_6144[4726] = ci_6144[698];
	assign cj_6144[4727] = ci_6144[4129];
	assign cj_6144[4728] = ci_6144[2376];
	assign cj_6144[4729] = ci_6144[1583];
	assign cj_6144[4730] = ci_6144[1750];
	assign cj_6144[4731] = ci_6144[2877];
	assign cj_6144[4732] = ci_6144[4964];
	assign cj_6144[4733] = ci_6144[1867];
	assign cj_6144[4734] = ci_6144[5874];
	assign cj_6144[4735] = ci_6144[4697];
	assign cj_6144[4736] = ci_6144[4480];
	assign cj_6144[4737] = ci_6144[5223];
	assign cj_6144[4738] = ci_6144[782];
	assign cj_6144[4739] = ci_6144[3445];
	assign cj_6144[4740] = ci_6144[924];
	assign cj_6144[4741] = ci_6144[5507];
	assign cj_6144[4742] = ci_6144[4906];
	assign cj_6144[4743] = ci_6144[5265];
	assign cj_6144[4744] = ci_6144[440];
	assign cj_6144[4745] = ci_6144[2719];
	assign cj_6144[4746] = ci_6144[5958];
	assign cj_6144[4747] = ci_6144[4013];
	assign cj_6144[4748] = ci_6144[3028];
	assign cj_6144[4749] = ci_6144[3003];
	assign cj_6144[4750] = ci_6144[3938];
	assign cj_6144[4751] = ci_6144[5833];
	assign cj_6144[4752] = ci_6144[2544];
	assign cj_6144[4753] = ci_6144[215];
	assign cj_6144[4754] = ci_6144[4990];
	assign cj_6144[4755] = ci_6144[4581];
	assign cj_6144[4756] = ci_6144[5132];
	assign cj_6144[4757] = ci_6144[499];
	assign cj_6144[4758] = ci_6144[2970];
	assign cj_6144[4759] = ci_6144[257];
	assign cj_6144[4760] = ci_6144[4648];
	assign cj_6144[4761] = ci_6144[3855];
	assign cj_6144[4762] = ci_6144[4022];
	assign cj_6144[4763] = ci_6144[5149];
	assign cj_6144[4764] = ci_6144[1092];
	assign cj_6144[4765] = ci_6144[4139];
	assign cj_6144[4766] = ci_6144[2002];
	assign cj_6144[4767] = ci_6144[825];
	assign cj_6144[4768] = ci_6144[608];
	assign cj_6144[4769] = ci_6144[1351];
	assign cj_6144[4770] = ci_6144[3054];
	assign cj_6144[4771] = ci_6144[5717];
	assign cj_6144[4772] = ci_6144[3196];
	assign cj_6144[4773] = ci_6144[1635];
	assign cj_6144[4774] = ci_6144[1034];
	assign cj_6144[4775] = ci_6144[1393];
	assign cj_6144[4776] = ci_6144[2712];
	assign cj_6144[4777] = ci_6144[4991];
	assign cj_6144[4778] = ci_6144[2086];
	assign cj_6144[4779] = ci_6144[141];
	assign cj_6144[4780] = ci_6144[5300];
	assign cj_6144[4781] = ci_6144[5275];
	assign cj_6144[4782] = ci_6144[66];
	assign cj_6144[4783] = ci_6144[1961];
	assign cj_6144[4784] = ci_6144[4816];
	assign cj_6144[4785] = ci_6144[2487];
	assign cj_6144[4786] = ci_6144[1118];
	assign cj_6144[4787] = ci_6144[709];
	assign cj_6144[4788] = ci_6144[1260];
	assign cj_6144[4789] = ci_6144[2771];
	assign cj_6144[4790] = ci_6144[5242];
	assign cj_6144[4791] = ci_6144[2529];
	assign cj_6144[4792] = ci_6144[776];
	assign cj_6144[4793] = ci_6144[6127];
	assign cj_6144[4794] = ci_6144[150];
	assign cj_6144[4795] = ci_6144[1277];
	assign cj_6144[4796] = ci_6144[3364];
	assign cj_6144[4797] = ci_6144[267];
	assign cj_6144[4798] = ci_6144[4274];
	assign cj_6144[4799] = ci_6144[3097];
	assign cj_6144[4800] = ci_6144[2880];
	assign cj_6144[4801] = ci_6144[3623];
	assign cj_6144[4802] = ci_6144[5326];
	assign cj_6144[4803] = ci_6144[1845];
	assign cj_6144[4804] = ci_6144[5468];
	assign cj_6144[4805] = ci_6144[3907];
	assign cj_6144[4806] = ci_6144[3306];
	assign cj_6144[4807] = ci_6144[3665];
	assign cj_6144[4808] = ci_6144[4984];
	assign cj_6144[4809] = ci_6144[1119];
	assign cj_6144[4810] = ci_6144[4358];
	assign cj_6144[4811] = ci_6144[2413];
	assign cj_6144[4812] = ci_6144[1428];
	assign cj_6144[4813] = ci_6144[1403];
	assign cj_6144[4814] = ci_6144[2338];
	assign cj_6144[4815] = ci_6144[4233];
	assign cj_6144[4816] = ci_6144[944];
	assign cj_6144[4817] = ci_6144[4759];
	assign cj_6144[4818] = ci_6144[3390];
	assign cj_6144[4819] = ci_6144[2981];
	assign cj_6144[4820] = ci_6144[3532];
	assign cj_6144[4821] = ci_6144[5043];
	assign cj_6144[4822] = ci_6144[1370];
	assign cj_6144[4823] = ci_6144[4801];
	assign cj_6144[4824] = ci_6144[3048];
	assign cj_6144[4825] = ci_6144[2255];
	assign cj_6144[4826] = ci_6144[2422];
	assign cj_6144[4827] = ci_6144[3549];
	assign cj_6144[4828] = ci_6144[5636];
	assign cj_6144[4829] = ci_6144[2539];
	assign cj_6144[4830] = ci_6144[402];
	assign cj_6144[4831] = ci_6144[5369];
	assign cj_6144[4832] = ci_6144[5152];
	assign cj_6144[4833] = ci_6144[5895];
	assign cj_6144[4834] = ci_6144[1454];
	assign cj_6144[4835] = ci_6144[4117];
	assign cj_6144[4836] = ci_6144[1596];
	assign cj_6144[4837] = ci_6144[35];
	assign cj_6144[4838] = ci_6144[5578];
	assign cj_6144[4839] = ci_6144[5937];
	assign cj_6144[4840] = ci_6144[1112];
	assign cj_6144[4841] = ci_6144[3391];
	assign cj_6144[4842] = ci_6144[486];
	assign cj_6144[4843] = ci_6144[4685];
	assign cj_6144[4844] = ci_6144[3700];
	assign cj_6144[4845] = ci_6144[3675];
	assign cj_6144[4846] = ci_6144[4610];
	assign cj_6144[4847] = ci_6144[361];
	assign cj_6144[4848] = ci_6144[3216];
	assign cj_6144[4849] = ci_6144[887];
	assign cj_6144[4850] = ci_6144[5662];
	assign cj_6144[4851] = ci_6144[5253];
	assign cj_6144[4852] = ci_6144[5804];
	assign cj_6144[4853] = ci_6144[1171];
	assign cj_6144[4854] = ci_6144[3642];
	assign cj_6144[4855] = ci_6144[929];
	assign cj_6144[4856] = ci_6144[5320];
	assign cj_6144[4857] = ci_6144[4527];
	assign cj_6144[4858] = ci_6144[4694];
	assign cj_6144[4859] = ci_6144[5821];
	assign cj_6144[4860] = ci_6144[1764];
	assign cj_6144[4861] = ci_6144[4811];
	assign cj_6144[4862] = ci_6144[2674];
	assign cj_6144[4863] = ci_6144[1497];
	assign cj_6144[4864] = ci_6144[1280];
	assign cj_6144[4865] = ci_6144[2023];
	assign cj_6144[4866] = ci_6144[3726];
	assign cj_6144[4867] = ci_6144[245];
	assign cj_6144[4868] = ci_6144[3868];
	assign cj_6144[4869] = ci_6144[2307];
	assign cj_6144[4870] = ci_6144[1706];
	assign cj_6144[4871] = ci_6144[2065];
	assign cj_6144[4872] = ci_6144[3384];
	assign cj_6144[4873] = ci_6144[5663];
	assign cj_6144[4874] = ci_6144[2758];
	assign cj_6144[4875] = ci_6144[813];
	assign cj_6144[4876] = ci_6144[5972];
	assign cj_6144[4877] = ci_6144[5947];
	assign cj_6144[4878] = ci_6144[738];
	assign cj_6144[4879] = ci_6144[2633];
	assign cj_6144[4880] = ci_6144[5488];
	assign cj_6144[4881] = ci_6144[3159];
	assign cj_6144[4882] = ci_6144[1790];
	assign cj_6144[4883] = ci_6144[1381];
	assign cj_6144[4884] = ci_6144[1932];
	assign cj_6144[4885] = ci_6144[3443];
	assign cj_6144[4886] = ci_6144[5914];
	assign cj_6144[4887] = ci_6144[3201];
	assign cj_6144[4888] = ci_6144[1448];
	assign cj_6144[4889] = ci_6144[655];
	assign cj_6144[4890] = ci_6144[822];
	assign cj_6144[4891] = ci_6144[1949];
	assign cj_6144[4892] = ci_6144[4036];
	assign cj_6144[4893] = ci_6144[939];
	assign cj_6144[4894] = ci_6144[4946];
	assign cj_6144[4895] = ci_6144[3769];
	assign cj_6144[4896] = ci_6144[3552];
	assign cj_6144[4897] = ci_6144[4295];
	assign cj_6144[4898] = ci_6144[5998];
	assign cj_6144[4899] = ci_6144[2517];
	assign cj_6144[4900] = ci_6144[6140];
	assign cj_6144[4901] = ci_6144[4579];
	assign cj_6144[4902] = ci_6144[3978];
	assign cj_6144[4903] = ci_6144[4337];
	assign cj_6144[4904] = ci_6144[5656];
	assign cj_6144[4905] = ci_6144[1791];
	assign cj_6144[4906] = ci_6144[5030];
	assign cj_6144[4907] = ci_6144[3085];
	assign cj_6144[4908] = ci_6144[2100];
	assign cj_6144[4909] = ci_6144[2075];
	assign cj_6144[4910] = ci_6144[3010];
	assign cj_6144[4911] = ci_6144[4905];
	assign cj_6144[4912] = ci_6144[1616];
	assign cj_6144[4913] = ci_6144[5431];
	assign cj_6144[4914] = ci_6144[4062];
	assign cj_6144[4915] = ci_6144[3653];
	assign cj_6144[4916] = ci_6144[4204];
	assign cj_6144[4917] = ci_6144[5715];
	assign cj_6144[4918] = ci_6144[2042];
	assign cj_6144[4919] = ci_6144[5473];
	assign cj_6144[4920] = ci_6144[3720];
	assign cj_6144[4921] = ci_6144[2927];
	assign cj_6144[4922] = ci_6144[3094];
	assign cj_6144[4923] = ci_6144[4221];
	assign cj_6144[4924] = ci_6144[164];
	assign cj_6144[4925] = ci_6144[3211];
	assign cj_6144[4926] = ci_6144[1074];
	assign cj_6144[4927] = ci_6144[6041];
	assign cj_6144[4928] = ci_6144[5824];
	assign cj_6144[4929] = ci_6144[423];
	assign cj_6144[4930] = ci_6144[2126];
	assign cj_6144[4931] = ci_6144[4789];
	assign cj_6144[4932] = ci_6144[2268];
	assign cj_6144[4933] = ci_6144[707];
	assign cj_6144[4934] = ci_6144[106];
	assign cj_6144[4935] = ci_6144[465];
	assign cj_6144[4936] = ci_6144[1784];
	assign cj_6144[4937] = ci_6144[4063];
	assign cj_6144[4938] = ci_6144[1158];
	assign cj_6144[4939] = ci_6144[5357];
	assign cj_6144[4940] = ci_6144[4372];
	assign cj_6144[4941] = ci_6144[4347];
	assign cj_6144[4942] = ci_6144[5282];
	assign cj_6144[4943] = ci_6144[1033];
	assign cj_6144[4944] = ci_6144[3888];
	assign cj_6144[4945] = ci_6144[1559];
	assign cj_6144[4946] = ci_6144[190];
	assign cj_6144[4947] = ci_6144[5925];
	assign cj_6144[4948] = ci_6144[332];
	assign cj_6144[4949] = ci_6144[1843];
	assign cj_6144[4950] = ci_6144[4314];
	assign cj_6144[4951] = ci_6144[1601];
	assign cj_6144[4952] = ci_6144[5992];
	assign cj_6144[4953] = ci_6144[5199];
	assign cj_6144[4954] = ci_6144[5366];
	assign cj_6144[4955] = ci_6144[349];
	assign cj_6144[4956] = ci_6144[2436];
	assign cj_6144[4957] = ci_6144[5483];
	assign cj_6144[4958] = ci_6144[3346];
	assign cj_6144[4959] = ci_6144[2169];
	assign cj_6144[4960] = ci_6144[1952];
	assign cj_6144[4961] = ci_6144[2695];
	assign cj_6144[4962] = ci_6144[4398];
	assign cj_6144[4963] = ci_6144[917];
	assign cj_6144[4964] = ci_6144[4540];
	assign cj_6144[4965] = ci_6144[2979];
	assign cj_6144[4966] = ci_6144[2378];
	assign cj_6144[4967] = ci_6144[2737];
	assign cj_6144[4968] = ci_6144[4056];
	assign cj_6144[4969] = ci_6144[191];
	assign cj_6144[4970] = ci_6144[3430];
	assign cj_6144[4971] = ci_6144[1485];
	assign cj_6144[4972] = ci_6144[500];
	assign cj_6144[4973] = ci_6144[475];
	assign cj_6144[4974] = ci_6144[1410];
	assign cj_6144[4975] = ci_6144[3305];
	assign cj_6144[4976] = ci_6144[16];
	assign cj_6144[4977] = ci_6144[3831];
	assign cj_6144[4978] = ci_6144[2462];
	assign cj_6144[4979] = ci_6144[2053];
	assign cj_6144[4980] = ci_6144[2604];
	assign cj_6144[4981] = ci_6144[4115];
	assign cj_6144[4982] = ci_6144[442];
	assign cj_6144[4983] = ci_6144[3873];
	assign cj_6144[4984] = ci_6144[2120];
	assign cj_6144[4985] = ci_6144[1327];
	assign cj_6144[4986] = ci_6144[1494];
	assign cj_6144[4987] = ci_6144[2621];
	assign cj_6144[4988] = ci_6144[4708];
	assign cj_6144[4989] = ci_6144[1611];
	assign cj_6144[4990] = ci_6144[5618];
	assign cj_6144[4991] = ci_6144[4441];
	assign cj_6144[4992] = ci_6144[4224];
	assign cj_6144[4993] = ci_6144[4967];
	assign cj_6144[4994] = ci_6144[526];
	assign cj_6144[4995] = ci_6144[3189];
	assign cj_6144[4996] = ci_6144[668];
	assign cj_6144[4997] = ci_6144[5251];
	assign cj_6144[4998] = ci_6144[4650];
	assign cj_6144[4999] = ci_6144[5009];
	assign cj_6144[5000] = ci_6144[184];
	assign cj_6144[5001] = ci_6144[2463];
	assign cj_6144[5002] = ci_6144[5702];
	assign cj_6144[5003] = ci_6144[3757];
	assign cj_6144[5004] = ci_6144[2772];
	assign cj_6144[5005] = ci_6144[2747];
	assign cj_6144[5006] = ci_6144[3682];
	assign cj_6144[5007] = ci_6144[5577];
	assign cj_6144[5008] = ci_6144[2288];
	assign cj_6144[5009] = ci_6144[6103];
	assign cj_6144[5010] = ci_6144[4734];
	assign cj_6144[5011] = ci_6144[4325];
	assign cj_6144[5012] = ci_6144[4876];
	assign cj_6144[5013] = ci_6144[243];
	assign cj_6144[5014] = ci_6144[2714];
	assign cj_6144[5015] = ci_6144[1];
	assign cj_6144[5016] = ci_6144[4392];
	assign cj_6144[5017] = ci_6144[3599];
	assign cj_6144[5018] = ci_6144[3766];
	assign cj_6144[5019] = ci_6144[4893];
	assign cj_6144[5020] = ci_6144[836];
	assign cj_6144[5021] = ci_6144[3883];
	assign cj_6144[5022] = ci_6144[1746];
	assign cj_6144[5023] = ci_6144[569];
	assign cj_6144[5024] = ci_6144[352];
	assign cj_6144[5025] = ci_6144[1095];
	assign cj_6144[5026] = ci_6144[2798];
	assign cj_6144[5027] = ci_6144[5461];
	assign cj_6144[5028] = ci_6144[2940];
	assign cj_6144[5029] = ci_6144[1379];
	assign cj_6144[5030] = ci_6144[778];
	assign cj_6144[5031] = ci_6144[1137];
	assign cj_6144[5032] = ci_6144[2456];
	assign cj_6144[5033] = ci_6144[4735];
	assign cj_6144[5034] = ci_6144[1830];
	assign cj_6144[5035] = ci_6144[6029];
	assign cj_6144[5036] = ci_6144[5044];
	assign cj_6144[5037] = ci_6144[5019];
	assign cj_6144[5038] = ci_6144[5954];
	assign cj_6144[5039] = ci_6144[1705];
	assign cj_6144[5040] = ci_6144[4560];
	assign cj_6144[5041] = ci_6144[2231];
	assign cj_6144[5042] = ci_6144[862];
	assign cj_6144[5043] = ci_6144[453];
	assign cj_6144[5044] = ci_6144[1004];
	assign cj_6144[5045] = ci_6144[2515];
	assign cj_6144[5046] = ci_6144[4986];
	assign cj_6144[5047] = ci_6144[2273];
	assign cj_6144[5048] = ci_6144[520];
	assign cj_6144[5049] = ci_6144[5871];
	assign cj_6144[5050] = ci_6144[6038];
	assign cj_6144[5051] = ci_6144[1021];
	assign cj_6144[5052] = ci_6144[3108];
	assign cj_6144[5053] = ci_6144[11];
	assign cj_6144[5054] = ci_6144[4018];
	assign cj_6144[5055] = ci_6144[2841];
	assign cj_6144[5056] = ci_6144[2624];
	assign cj_6144[5057] = ci_6144[3367];
	assign cj_6144[5058] = ci_6144[5070];
	assign cj_6144[5059] = ci_6144[1589];
	assign cj_6144[5060] = ci_6144[5212];
	assign cj_6144[5061] = ci_6144[3651];
	assign cj_6144[5062] = ci_6144[3050];
	assign cj_6144[5063] = ci_6144[3409];
	assign cj_6144[5064] = ci_6144[4728];
	assign cj_6144[5065] = ci_6144[863];
	assign cj_6144[5066] = ci_6144[4102];
	assign cj_6144[5067] = ci_6144[2157];
	assign cj_6144[5068] = ci_6144[1172];
	assign cj_6144[5069] = ci_6144[1147];
	assign cj_6144[5070] = ci_6144[2082];
	assign cj_6144[5071] = ci_6144[3977];
	assign cj_6144[5072] = ci_6144[688];
	assign cj_6144[5073] = ci_6144[4503];
	assign cj_6144[5074] = ci_6144[3134];
	assign cj_6144[5075] = ci_6144[2725];
	assign cj_6144[5076] = ci_6144[3276];
	assign cj_6144[5077] = ci_6144[4787];
	assign cj_6144[5078] = ci_6144[1114];
	assign cj_6144[5079] = ci_6144[4545];
	assign cj_6144[5080] = ci_6144[2792];
	assign cj_6144[5081] = ci_6144[1999];
	assign cj_6144[5082] = ci_6144[2166];
	assign cj_6144[5083] = ci_6144[3293];
	assign cj_6144[5084] = ci_6144[5380];
	assign cj_6144[5085] = ci_6144[2283];
	assign cj_6144[5086] = ci_6144[146];
	assign cj_6144[5087] = ci_6144[5113];
	assign cj_6144[5088] = ci_6144[4896];
	assign cj_6144[5089] = ci_6144[5639];
	assign cj_6144[5090] = ci_6144[1198];
	assign cj_6144[5091] = ci_6144[3861];
	assign cj_6144[5092] = ci_6144[1340];
	assign cj_6144[5093] = ci_6144[5923];
	assign cj_6144[5094] = ci_6144[5322];
	assign cj_6144[5095] = ci_6144[5681];
	assign cj_6144[5096] = ci_6144[856];
	assign cj_6144[5097] = ci_6144[3135];
	assign cj_6144[5098] = ci_6144[230];
	assign cj_6144[5099] = ci_6144[4429];
	assign cj_6144[5100] = ci_6144[3444];
	assign cj_6144[5101] = ci_6144[3419];
	assign cj_6144[5102] = ci_6144[4354];
	assign cj_6144[5103] = ci_6144[105];
	assign cj_6144[5104] = ci_6144[2960];
	assign cj_6144[5105] = ci_6144[631];
	assign cj_6144[5106] = ci_6144[5406];
	assign cj_6144[5107] = ci_6144[4997];
	assign cj_6144[5108] = ci_6144[5548];
	assign cj_6144[5109] = ci_6144[915];
	assign cj_6144[5110] = ci_6144[3386];
	assign cj_6144[5111] = ci_6144[673];
	assign cj_6144[5112] = ci_6144[5064];
	assign cj_6144[5113] = ci_6144[4271];
	assign cj_6144[5114] = ci_6144[4438];
	assign cj_6144[5115] = ci_6144[5565];
	assign cj_6144[5116] = ci_6144[1508];
	assign cj_6144[5117] = ci_6144[4555];
	assign cj_6144[5118] = ci_6144[2418];
	assign cj_6144[5119] = ci_6144[1241];
	assign cj_6144[5120] = ci_6144[1024];
	assign cj_6144[5121] = ci_6144[1767];
	assign cj_6144[5122] = ci_6144[3470];
	assign cj_6144[5123] = ci_6144[6133];
	assign cj_6144[5124] = ci_6144[3612];
	assign cj_6144[5125] = ci_6144[2051];
	assign cj_6144[5126] = ci_6144[1450];
	assign cj_6144[5127] = ci_6144[1809];
	assign cj_6144[5128] = ci_6144[3128];
	assign cj_6144[5129] = ci_6144[5407];
	assign cj_6144[5130] = ci_6144[2502];
	assign cj_6144[5131] = ci_6144[557];
	assign cj_6144[5132] = ci_6144[5716];
	assign cj_6144[5133] = ci_6144[5691];
	assign cj_6144[5134] = ci_6144[482];
	assign cj_6144[5135] = ci_6144[2377];
	assign cj_6144[5136] = ci_6144[5232];
	assign cj_6144[5137] = ci_6144[2903];
	assign cj_6144[5138] = ci_6144[1534];
	assign cj_6144[5139] = ci_6144[1125];
	assign cj_6144[5140] = ci_6144[1676];
	assign cj_6144[5141] = ci_6144[3187];
	assign cj_6144[5142] = ci_6144[5658];
	assign cj_6144[5143] = ci_6144[2945];
	assign cj_6144[5144] = ci_6144[1192];
	assign cj_6144[5145] = ci_6144[399];
	assign cj_6144[5146] = ci_6144[566];
	assign cj_6144[5147] = ci_6144[1693];
	assign cj_6144[5148] = ci_6144[3780];
	assign cj_6144[5149] = ci_6144[683];
	assign cj_6144[5150] = ci_6144[4690];
	assign cj_6144[5151] = ci_6144[3513];
	assign cj_6144[5152] = ci_6144[3296];
	assign cj_6144[5153] = ci_6144[4039];
	assign cj_6144[5154] = ci_6144[5742];
	assign cj_6144[5155] = ci_6144[2261];
	assign cj_6144[5156] = ci_6144[5884];
	assign cj_6144[5157] = ci_6144[4323];
	assign cj_6144[5158] = ci_6144[3722];
	assign cj_6144[5159] = ci_6144[4081];
	assign cj_6144[5160] = ci_6144[5400];
	assign cj_6144[5161] = ci_6144[1535];
	assign cj_6144[5162] = ci_6144[4774];
	assign cj_6144[5163] = ci_6144[2829];
	assign cj_6144[5164] = ci_6144[1844];
	assign cj_6144[5165] = ci_6144[1819];
	assign cj_6144[5166] = ci_6144[2754];
	assign cj_6144[5167] = ci_6144[4649];
	assign cj_6144[5168] = ci_6144[1360];
	assign cj_6144[5169] = ci_6144[5175];
	assign cj_6144[5170] = ci_6144[3806];
	assign cj_6144[5171] = ci_6144[3397];
	assign cj_6144[5172] = ci_6144[3948];
	assign cj_6144[5173] = ci_6144[5459];
	assign cj_6144[5174] = ci_6144[1786];
	assign cj_6144[5175] = ci_6144[5217];
	assign cj_6144[5176] = ci_6144[3464];
	assign cj_6144[5177] = ci_6144[2671];
	assign cj_6144[5178] = ci_6144[2838];
	assign cj_6144[5179] = ci_6144[3965];
	assign cj_6144[5180] = ci_6144[6052];
	assign cj_6144[5181] = ci_6144[2955];
	assign cj_6144[5182] = ci_6144[818];
	assign cj_6144[5183] = ci_6144[5785];
	assign cj_6144[5184] = ci_6144[5568];
	assign cj_6144[5185] = ci_6144[167];
	assign cj_6144[5186] = ci_6144[1870];
	assign cj_6144[5187] = ci_6144[4533];
	assign cj_6144[5188] = ci_6144[2012];
	assign cj_6144[5189] = ci_6144[451];
	assign cj_6144[5190] = ci_6144[5994];
	assign cj_6144[5191] = ci_6144[209];
	assign cj_6144[5192] = ci_6144[1528];
	assign cj_6144[5193] = ci_6144[3807];
	assign cj_6144[5194] = ci_6144[902];
	assign cj_6144[5195] = ci_6144[5101];
	assign cj_6144[5196] = ci_6144[4116];
	assign cj_6144[5197] = ci_6144[4091];
	assign cj_6144[5198] = ci_6144[5026];
	assign cj_6144[5199] = ci_6144[777];
	assign cj_6144[5200] = ci_6144[3632];
	assign cj_6144[5201] = ci_6144[1303];
	assign cj_6144[5202] = ci_6144[6078];
	assign cj_6144[5203] = ci_6144[5669];
	assign cj_6144[5204] = ci_6144[76];
	assign cj_6144[5205] = ci_6144[1587];
	assign cj_6144[5206] = ci_6144[4058];
	assign cj_6144[5207] = ci_6144[1345];
	assign cj_6144[5208] = ci_6144[5736];
	assign cj_6144[5209] = ci_6144[4943];
	assign cj_6144[5210] = ci_6144[5110];
	assign cj_6144[5211] = ci_6144[93];
	assign cj_6144[5212] = ci_6144[2180];
	assign cj_6144[5213] = ci_6144[5227];
	assign cj_6144[5214] = ci_6144[3090];
	assign cj_6144[5215] = ci_6144[1913];
	assign cj_6144[5216] = ci_6144[1696];
	assign cj_6144[5217] = ci_6144[2439];
	assign cj_6144[5218] = ci_6144[4142];
	assign cj_6144[5219] = ci_6144[661];
	assign cj_6144[5220] = ci_6144[4284];
	assign cj_6144[5221] = ci_6144[2723];
	assign cj_6144[5222] = ci_6144[2122];
	assign cj_6144[5223] = ci_6144[2481];
	assign cj_6144[5224] = ci_6144[3800];
	assign cj_6144[5225] = ci_6144[6079];
	assign cj_6144[5226] = ci_6144[3174];
	assign cj_6144[5227] = ci_6144[1229];
	assign cj_6144[5228] = ci_6144[244];
	assign cj_6144[5229] = ci_6144[219];
	assign cj_6144[5230] = ci_6144[1154];
	assign cj_6144[5231] = ci_6144[3049];
	assign cj_6144[5232] = ci_6144[5904];
	assign cj_6144[5233] = ci_6144[3575];
	assign cj_6144[5234] = ci_6144[2206];
	assign cj_6144[5235] = ci_6144[1797];
	assign cj_6144[5236] = ci_6144[2348];
	assign cj_6144[5237] = ci_6144[3859];
	assign cj_6144[5238] = ci_6144[186];
	assign cj_6144[5239] = ci_6144[3617];
	assign cj_6144[5240] = ci_6144[1864];
	assign cj_6144[5241] = ci_6144[1071];
	assign cj_6144[5242] = ci_6144[1238];
	assign cj_6144[5243] = ci_6144[2365];
	assign cj_6144[5244] = ci_6144[4452];
	assign cj_6144[5245] = ci_6144[1355];
	assign cj_6144[5246] = ci_6144[5362];
	assign cj_6144[5247] = ci_6144[4185];
	assign cj_6144[5248] = ci_6144[3968];
	assign cj_6144[5249] = ci_6144[4711];
	assign cj_6144[5250] = ci_6144[270];
	assign cj_6144[5251] = ci_6144[2933];
	assign cj_6144[5252] = ci_6144[412];
	assign cj_6144[5253] = ci_6144[4995];
	assign cj_6144[5254] = ci_6144[4394];
	assign cj_6144[5255] = ci_6144[4753];
	assign cj_6144[5256] = ci_6144[6072];
	assign cj_6144[5257] = ci_6144[2207];
	assign cj_6144[5258] = ci_6144[5446];
	assign cj_6144[5259] = ci_6144[3501];
	assign cj_6144[5260] = ci_6144[2516];
	assign cj_6144[5261] = ci_6144[2491];
	assign cj_6144[5262] = ci_6144[3426];
	assign cj_6144[5263] = ci_6144[5321];
	assign cj_6144[5264] = ci_6144[2032];
	assign cj_6144[5265] = ci_6144[5847];
	assign cj_6144[5266] = ci_6144[4478];
	assign cj_6144[5267] = ci_6144[4069];
	assign cj_6144[5268] = ci_6144[4620];
	assign cj_6144[5269] = ci_6144[6131];
	assign cj_6144[5270] = ci_6144[2458];
	assign cj_6144[5271] = ci_6144[5889];
	assign cj_6144[5272] = ci_6144[4136];
	assign cj_6144[5273] = ci_6144[3343];
	assign cj_6144[5274] = ci_6144[3510];
	assign cj_6144[5275] = ci_6144[4637];
	assign cj_6144[5276] = ci_6144[580];
	assign cj_6144[5277] = ci_6144[3627];
	assign cj_6144[5278] = ci_6144[1490];
	assign cj_6144[5279] = ci_6144[313];
	assign cj_6144[5280] = ci_6144[96];
	assign cj_6144[5281] = ci_6144[839];
	assign cj_6144[5282] = ci_6144[2542];
	assign cj_6144[5283] = ci_6144[5205];
	assign cj_6144[5284] = ci_6144[2684];
	assign cj_6144[5285] = ci_6144[1123];
	assign cj_6144[5286] = ci_6144[522];
	assign cj_6144[5287] = ci_6144[881];
	assign cj_6144[5288] = ci_6144[2200];
	assign cj_6144[5289] = ci_6144[4479];
	assign cj_6144[5290] = ci_6144[1574];
	assign cj_6144[5291] = ci_6144[5773];
	assign cj_6144[5292] = ci_6144[4788];
	assign cj_6144[5293] = ci_6144[4763];
	assign cj_6144[5294] = ci_6144[5698];
	assign cj_6144[5295] = ci_6144[1449];
	assign cj_6144[5296] = ci_6144[4304];
	assign cj_6144[5297] = ci_6144[1975];
	assign cj_6144[5298] = ci_6144[606];
	assign cj_6144[5299] = ci_6144[197];
	assign cj_6144[5300] = ci_6144[748];
	assign cj_6144[5301] = ci_6144[2259];
	assign cj_6144[5302] = ci_6144[4730];
	assign cj_6144[5303] = ci_6144[2017];
	assign cj_6144[5304] = ci_6144[264];
	assign cj_6144[5305] = ci_6144[5615];
	assign cj_6144[5306] = ci_6144[5782];
	assign cj_6144[5307] = ci_6144[765];
	assign cj_6144[5308] = ci_6144[2852];
	assign cj_6144[5309] = ci_6144[5899];
	assign cj_6144[5310] = ci_6144[3762];
	assign cj_6144[5311] = ci_6144[2585];
	assign cj_6144[5312] = ci_6144[2368];
	assign cj_6144[5313] = ci_6144[3111];
	assign cj_6144[5314] = ci_6144[4814];
	assign cj_6144[5315] = ci_6144[1333];
	assign cj_6144[5316] = ci_6144[4956];
	assign cj_6144[5317] = ci_6144[3395];
	assign cj_6144[5318] = ci_6144[2794];
	assign cj_6144[5319] = ci_6144[3153];
	assign cj_6144[5320] = ci_6144[4472];
	assign cj_6144[5321] = ci_6144[607];
	assign cj_6144[5322] = ci_6144[3846];
	assign cj_6144[5323] = ci_6144[1901];
	assign cj_6144[5324] = ci_6144[916];
	assign cj_6144[5325] = ci_6144[891];
	assign cj_6144[5326] = ci_6144[1826];
	assign cj_6144[5327] = ci_6144[3721];
	assign cj_6144[5328] = ci_6144[432];
	assign cj_6144[5329] = ci_6144[4247];
	assign cj_6144[5330] = ci_6144[2878];
	assign cj_6144[5331] = ci_6144[2469];
	assign cj_6144[5332] = ci_6144[3020];
	assign cj_6144[5333] = ci_6144[4531];
	assign cj_6144[5334] = ci_6144[858];
	assign cj_6144[5335] = ci_6144[4289];
	assign cj_6144[5336] = ci_6144[2536];
	assign cj_6144[5337] = ci_6144[1743];
	assign cj_6144[5338] = ci_6144[1910];
	assign cj_6144[5339] = ci_6144[3037];
	assign cj_6144[5340] = ci_6144[5124];
	assign cj_6144[5341] = ci_6144[2027];
	assign cj_6144[5342] = ci_6144[6034];
	assign cj_6144[5343] = ci_6144[4857];
	assign cj_6144[5344] = ci_6144[4640];
	assign cj_6144[5345] = ci_6144[5383];
	assign cj_6144[5346] = ci_6144[942];
	assign cj_6144[5347] = ci_6144[3605];
	assign cj_6144[5348] = ci_6144[1084];
	assign cj_6144[5349] = ci_6144[5667];
	assign cj_6144[5350] = ci_6144[5066];
	assign cj_6144[5351] = ci_6144[5425];
	assign cj_6144[5352] = ci_6144[600];
	assign cj_6144[5353] = ci_6144[2879];
	assign cj_6144[5354] = ci_6144[6118];
	assign cj_6144[5355] = ci_6144[4173];
	assign cj_6144[5356] = ci_6144[3188];
	assign cj_6144[5357] = ci_6144[3163];
	assign cj_6144[5358] = ci_6144[4098];
	assign cj_6144[5359] = ci_6144[5993];
	assign cj_6144[5360] = ci_6144[2704];
	assign cj_6144[5361] = ci_6144[375];
	assign cj_6144[5362] = ci_6144[5150];
	assign cj_6144[5363] = ci_6144[4741];
	assign cj_6144[5364] = ci_6144[5292];
	assign cj_6144[5365] = ci_6144[659];
	assign cj_6144[5366] = ci_6144[3130];
	assign cj_6144[5367] = ci_6144[417];
	assign cj_6144[5368] = ci_6144[4808];
	assign cj_6144[5369] = ci_6144[4015];
	assign cj_6144[5370] = ci_6144[4182];
	assign cj_6144[5371] = ci_6144[5309];
	assign cj_6144[5372] = ci_6144[1252];
	assign cj_6144[5373] = ci_6144[4299];
	assign cj_6144[5374] = ci_6144[2162];
	assign cj_6144[5375] = ci_6144[985];
	assign cj_6144[5376] = ci_6144[768];
	assign cj_6144[5377] = ci_6144[1511];
	assign cj_6144[5378] = ci_6144[3214];
	assign cj_6144[5379] = ci_6144[5877];
	assign cj_6144[5380] = ci_6144[3356];
	assign cj_6144[5381] = ci_6144[1795];
	assign cj_6144[5382] = ci_6144[1194];
	assign cj_6144[5383] = ci_6144[1553];
	assign cj_6144[5384] = ci_6144[2872];
	assign cj_6144[5385] = ci_6144[5151];
	assign cj_6144[5386] = ci_6144[2246];
	assign cj_6144[5387] = ci_6144[301];
	assign cj_6144[5388] = ci_6144[5460];
	assign cj_6144[5389] = ci_6144[5435];
	assign cj_6144[5390] = ci_6144[226];
	assign cj_6144[5391] = ci_6144[2121];
	assign cj_6144[5392] = ci_6144[4976];
	assign cj_6144[5393] = ci_6144[2647];
	assign cj_6144[5394] = ci_6144[1278];
	assign cj_6144[5395] = ci_6144[869];
	assign cj_6144[5396] = ci_6144[1420];
	assign cj_6144[5397] = ci_6144[2931];
	assign cj_6144[5398] = ci_6144[5402];
	assign cj_6144[5399] = ci_6144[2689];
	assign cj_6144[5400] = ci_6144[936];
	assign cj_6144[5401] = ci_6144[143];
	assign cj_6144[5402] = ci_6144[310];
	assign cj_6144[5403] = ci_6144[1437];
	assign cj_6144[5404] = ci_6144[3524];
	assign cj_6144[5405] = ci_6144[427];
	assign cj_6144[5406] = ci_6144[4434];
	assign cj_6144[5407] = ci_6144[3257];
	assign cj_6144[5408] = ci_6144[3040];
	assign cj_6144[5409] = ci_6144[3783];
	assign cj_6144[5410] = ci_6144[5486];
	assign cj_6144[5411] = ci_6144[2005];
	assign cj_6144[5412] = ci_6144[5628];
	assign cj_6144[5413] = ci_6144[4067];
	assign cj_6144[5414] = ci_6144[3466];
	assign cj_6144[5415] = ci_6144[3825];
	assign cj_6144[5416] = ci_6144[5144];
	assign cj_6144[5417] = ci_6144[1279];
	assign cj_6144[5418] = ci_6144[4518];
	assign cj_6144[5419] = ci_6144[2573];
	assign cj_6144[5420] = ci_6144[1588];
	assign cj_6144[5421] = ci_6144[1563];
	assign cj_6144[5422] = ci_6144[2498];
	assign cj_6144[5423] = ci_6144[4393];
	assign cj_6144[5424] = ci_6144[1104];
	assign cj_6144[5425] = ci_6144[4919];
	assign cj_6144[5426] = ci_6144[3550];
	assign cj_6144[5427] = ci_6144[3141];
	assign cj_6144[5428] = ci_6144[3692];
	assign cj_6144[5429] = ci_6144[5203];
	assign cj_6144[5430] = ci_6144[1530];
	assign cj_6144[5431] = ci_6144[4961];
	assign cj_6144[5432] = ci_6144[3208];
	assign cj_6144[5433] = ci_6144[2415];
	assign cj_6144[5434] = ci_6144[2582];
	assign cj_6144[5435] = ci_6144[3709];
	assign cj_6144[5436] = ci_6144[5796];
	assign cj_6144[5437] = ci_6144[2699];
	assign cj_6144[5438] = ci_6144[562];
	assign cj_6144[5439] = ci_6144[5529];
	assign cj_6144[5440] = ci_6144[5312];
	assign cj_6144[5441] = ci_6144[6055];
	assign cj_6144[5442] = ci_6144[1614];
	assign cj_6144[5443] = ci_6144[4277];
	assign cj_6144[5444] = ci_6144[1756];
	assign cj_6144[5445] = ci_6144[195];
	assign cj_6144[5446] = ci_6144[5738];
	assign cj_6144[5447] = ci_6144[6097];
	assign cj_6144[5448] = ci_6144[1272];
	assign cj_6144[5449] = ci_6144[3551];
	assign cj_6144[5450] = ci_6144[646];
	assign cj_6144[5451] = ci_6144[4845];
	assign cj_6144[5452] = ci_6144[3860];
	assign cj_6144[5453] = ci_6144[3835];
	assign cj_6144[5454] = ci_6144[4770];
	assign cj_6144[5455] = ci_6144[521];
	assign cj_6144[5456] = ci_6144[3376];
	assign cj_6144[5457] = ci_6144[1047];
	assign cj_6144[5458] = ci_6144[5822];
	assign cj_6144[5459] = ci_6144[5413];
	assign cj_6144[5460] = ci_6144[5964];
	assign cj_6144[5461] = ci_6144[1331];
	assign cj_6144[5462] = ci_6144[3802];
	assign cj_6144[5463] = ci_6144[1089];
	assign cj_6144[5464] = ci_6144[5480];
	assign cj_6144[5465] = ci_6144[4687];
	assign cj_6144[5466] = ci_6144[4854];
	assign cj_6144[5467] = ci_6144[5981];
	assign cj_6144[5468] = ci_6144[1924];
	assign cj_6144[5469] = ci_6144[4971];
	assign cj_6144[5470] = ci_6144[2834];
	assign cj_6144[5471] = ci_6144[1657];
	assign cj_6144[5472] = ci_6144[1440];
	assign cj_6144[5473] = ci_6144[2183];
	assign cj_6144[5474] = ci_6144[3886];
	assign cj_6144[5475] = ci_6144[405];
	assign cj_6144[5476] = ci_6144[4028];
	assign cj_6144[5477] = ci_6144[2467];
	assign cj_6144[5478] = ci_6144[1866];
	assign cj_6144[5479] = ci_6144[2225];
	assign cj_6144[5480] = ci_6144[3544];
	assign cj_6144[5481] = ci_6144[5823];
	assign cj_6144[5482] = ci_6144[2918];
	assign cj_6144[5483] = ci_6144[973];
	assign cj_6144[5484] = ci_6144[6132];
	assign cj_6144[5485] = ci_6144[6107];
	assign cj_6144[5486] = ci_6144[898];
	assign cj_6144[5487] = ci_6144[2793];
	assign cj_6144[5488] = ci_6144[5648];
	assign cj_6144[5489] = ci_6144[3319];
	assign cj_6144[5490] = ci_6144[1950];
	assign cj_6144[5491] = ci_6144[1541];
	assign cj_6144[5492] = ci_6144[2092];
	assign cj_6144[5493] = ci_6144[3603];
	assign cj_6144[5494] = ci_6144[6074];
	assign cj_6144[5495] = ci_6144[3361];
	assign cj_6144[5496] = ci_6144[1608];
	assign cj_6144[5497] = ci_6144[815];
	assign cj_6144[5498] = ci_6144[982];
	assign cj_6144[5499] = ci_6144[2109];
	assign cj_6144[5500] = ci_6144[4196];
	assign cj_6144[5501] = ci_6144[1099];
	assign cj_6144[5502] = ci_6144[5106];
	assign cj_6144[5503] = ci_6144[3929];
	assign cj_6144[5504] = ci_6144[3712];
	assign cj_6144[5505] = ci_6144[4455];
	assign cj_6144[5506] = ci_6144[14];
	assign cj_6144[5507] = ci_6144[2677];
	assign cj_6144[5508] = ci_6144[156];
	assign cj_6144[5509] = ci_6144[4739];
	assign cj_6144[5510] = ci_6144[4138];
	assign cj_6144[5511] = ci_6144[4497];
	assign cj_6144[5512] = ci_6144[5816];
	assign cj_6144[5513] = ci_6144[1951];
	assign cj_6144[5514] = ci_6144[5190];
	assign cj_6144[5515] = ci_6144[3245];
	assign cj_6144[5516] = ci_6144[2260];
	assign cj_6144[5517] = ci_6144[2235];
	assign cj_6144[5518] = ci_6144[3170];
	assign cj_6144[5519] = ci_6144[5065];
	assign cj_6144[5520] = ci_6144[1776];
	assign cj_6144[5521] = ci_6144[5591];
	assign cj_6144[5522] = ci_6144[4222];
	assign cj_6144[5523] = ci_6144[3813];
	assign cj_6144[5524] = ci_6144[4364];
	assign cj_6144[5525] = ci_6144[5875];
	assign cj_6144[5526] = ci_6144[2202];
	assign cj_6144[5527] = ci_6144[5633];
	assign cj_6144[5528] = ci_6144[3880];
	assign cj_6144[5529] = ci_6144[3087];
	assign cj_6144[5530] = ci_6144[3254];
	assign cj_6144[5531] = ci_6144[4381];
	assign cj_6144[5532] = ci_6144[324];
	assign cj_6144[5533] = ci_6144[3371];
	assign cj_6144[5534] = ci_6144[1234];
	assign cj_6144[5535] = ci_6144[57];
	assign cj_6144[5536] = ci_6144[5984];
	assign cj_6144[5537] = ci_6144[583];
	assign cj_6144[5538] = ci_6144[2286];
	assign cj_6144[5539] = ci_6144[4949];
	assign cj_6144[5540] = ci_6144[2428];
	assign cj_6144[5541] = ci_6144[867];
	assign cj_6144[5542] = ci_6144[266];
	assign cj_6144[5543] = ci_6144[625];
	assign cj_6144[5544] = ci_6144[1944];
	assign cj_6144[5545] = ci_6144[4223];
	assign cj_6144[5546] = ci_6144[1318];
	assign cj_6144[5547] = ci_6144[5517];
	assign cj_6144[5548] = ci_6144[4532];
	assign cj_6144[5549] = ci_6144[4507];
	assign cj_6144[5550] = ci_6144[5442];
	assign cj_6144[5551] = ci_6144[1193];
	assign cj_6144[5552] = ci_6144[4048];
	assign cj_6144[5553] = ci_6144[1719];
	assign cj_6144[5554] = ci_6144[350];
	assign cj_6144[5555] = ci_6144[6085];
	assign cj_6144[5556] = ci_6144[492];
	assign cj_6144[5557] = ci_6144[2003];
	assign cj_6144[5558] = ci_6144[4474];
	assign cj_6144[5559] = ci_6144[1761];
	assign cj_6144[5560] = ci_6144[8];
	assign cj_6144[5561] = ci_6144[5359];
	assign cj_6144[5562] = ci_6144[5526];
	assign cj_6144[5563] = ci_6144[509];
	assign cj_6144[5564] = ci_6144[2596];
	assign cj_6144[5565] = ci_6144[5643];
	assign cj_6144[5566] = ci_6144[3506];
	assign cj_6144[5567] = ci_6144[2329];
	assign cj_6144[5568] = ci_6144[2112];
	assign cj_6144[5569] = ci_6144[2855];
	assign cj_6144[5570] = ci_6144[4558];
	assign cj_6144[5571] = ci_6144[1077];
	assign cj_6144[5572] = ci_6144[4700];
	assign cj_6144[5573] = ci_6144[3139];
	assign cj_6144[5574] = ci_6144[2538];
	assign cj_6144[5575] = ci_6144[2897];
	assign cj_6144[5576] = ci_6144[4216];
	assign cj_6144[5577] = ci_6144[351];
	assign cj_6144[5578] = ci_6144[3590];
	assign cj_6144[5579] = ci_6144[1645];
	assign cj_6144[5580] = ci_6144[660];
	assign cj_6144[5581] = ci_6144[635];
	assign cj_6144[5582] = ci_6144[1570];
	assign cj_6144[5583] = ci_6144[3465];
	assign cj_6144[5584] = ci_6144[176];
	assign cj_6144[5585] = ci_6144[3991];
	assign cj_6144[5586] = ci_6144[2622];
	assign cj_6144[5587] = ci_6144[2213];
	assign cj_6144[5588] = ci_6144[2764];
	assign cj_6144[5589] = ci_6144[4275];
	assign cj_6144[5590] = ci_6144[602];
	assign cj_6144[5591] = ci_6144[4033];
	assign cj_6144[5592] = ci_6144[2280];
	assign cj_6144[5593] = ci_6144[1487];
	assign cj_6144[5594] = ci_6144[1654];
	assign cj_6144[5595] = ci_6144[2781];
	assign cj_6144[5596] = ci_6144[4868];
	assign cj_6144[5597] = ci_6144[1771];
	assign cj_6144[5598] = ci_6144[5778];
	assign cj_6144[5599] = ci_6144[4601];
	assign cj_6144[5600] = ci_6144[4384];
	assign cj_6144[5601] = ci_6144[5127];
	assign cj_6144[5602] = ci_6144[686];
	assign cj_6144[5603] = ci_6144[3349];
	assign cj_6144[5604] = ci_6144[828];
	assign cj_6144[5605] = ci_6144[5411];
	assign cj_6144[5606] = ci_6144[4810];
	assign cj_6144[5607] = ci_6144[5169];
	assign cj_6144[5608] = ci_6144[344];
	assign cj_6144[5609] = ci_6144[2623];
	assign cj_6144[5610] = ci_6144[5862];
	assign cj_6144[5611] = ci_6144[3917];
	assign cj_6144[5612] = ci_6144[2932];
	assign cj_6144[5613] = ci_6144[2907];
	assign cj_6144[5614] = ci_6144[3842];
	assign cj_6144[5615] = ci_6144[5737];
	assign cj_6144[5616] = ci_6144[2448];
	assign cj_6144[5617] = ci_6144[119];
	assign cj_6144[5618] = ci_6144[4894];
	assign cj_6144[5619] = ci_6144[4485];
	assign cj_6144[5620] = ci_6144[5036];
	assign cj_6144[5621] = ci_6144[403];
	assign cj_6144[5622] = ci_6144[2874];
	assign cj_6144[5623] = ci_6144[161];
	assign cj_6144[5624] = ci_6144[4552];
	assign cj_6144[5625] = ci_6144[3759];
	assign cj_6144[5626] = ci_6144[3926];
	assign cj_6144[5627] = ci_6144[5053];
	assign cj_6144[5628] = ci_6144[996];
	assign cj_6144[5629] = ci_6144[4043];
	assign cj_6144[5630] = ci_6144[1906];
	assign cj_6144[5631] = ci_6144[729];
	assign cj_6144[5632] = ci_6144[512];
	assign cj_6144[5633] = ci_6144[1255];
	assign cj_6144[5634] = ci_6144[2958];
	assign cj_6144[5635] = ci_6144[5621];
	assign cj_6144[5636] = ci_6144[3100];
	assign cj_6144[5637] = ci_6144[1539];
	assign cj_6144[5638] = ci_6144[938];
	assign cj_6144[5639] = ci_6144[1297];
	assign cj_6144[5640] = ci_6144[2616];
	assign cj_6144[5641] = ci_6144[4895];
	assign cj_6144[5642] = ci_6144[1990];
	assign cj_6144[5643] = ci_6144[45];
	assign cj_6144[5644] = ci_6144[5204];
	assign cj_6144[5645] = ci_6144[5179];
	assign cj_6144[5646] = ci_6144[6114];
	assign cj_6144[5647] = ci_6144[1865];
	assign cj_6144[5648] = ci_6144[4720];
	assign cj_6144[5649] = ci_6144[2391];
	assign cj_6144[5650] = ci_6144[1022];
	assign cj_6144[5651] = ci_6144[613];
	assign cj_6144[5652] = ci_6144[1164];
	assign cj_6144[5653] = ci_6144[2675];
	assign cj_6144[5654] = ci_6144[5146];
	assign cj_6144[5655] = ci_6144[2433];
	assign cj_6144[5656] = ci_6144[680];
	assign cj_6144[5657] = ci_6144[6031];
	assign cj_6144[5658] = ci_6144[54];
	assign cj_6144[5659] = ci_6144[1181];
	assign cj_6144[5660] = ci_6144[3268];
	assign cj_6144[5661] = ci_6144[171];
	assign cj_6144[5662] = ci_6144[4178];
	assign cj_6144[5663] = ci_6144[3001];
	assign cj_6144[5664] = ci_6144[2784];
	assign cj_6144[5665] = ci_6144[3527];
	assign cj_6144[5666] = ci_6144[5230];
	assign cj_6144[5667] = ci_6144[1749];
	assign cj_6144[5668] = ci_6144[5372];
	assign cj_6144[5669] = ci_6144[3811];
	assign cj_6144[5670] = ci_6144[3210];
	assign cj_6144[5671] = ci_6144[3569];
	assign cj_6144[5672] = ci_6144[4888];
	assign cj_6144[5673] = ci_6144[1023];
	assign cj_6144[5674] = ci_6144[4262];
	assign cj_6144[5675] = ci_6144[2317];
	assign cj_6144[5676] = ci_6144[1332];
	assign cj_6144[5677] = ci_6144[1307];
	assign cj_6144[5678] = ci_6144[2242];
	assign cj_6144[5679] = ci_6144[4137];
	assign cj_6144[5680] = ci_6144[848];
	assign cj_6144[5681] = ci_6144[4663];
	assign cj_6144[5682] = ci_6144[3294];
	assign cj_6144[5683] = ci_6144[2885];
	assign cj_6144[5684] = ci_6144[3436];
	assign cj_6144[5685] = ci_6144[4947];
	assign cj_6144[5686] = ci_6144[1274];
	assign cj_6144[5687] = ci_6144[4705];
	assign cj_6144[5688] = ci_6144[2952];
	assign cj_6144[5689] = ci_6144[2159];
	assign cj_6144[5690] = ci_6144[2326];
	assign cj_6144[5691] = ci_6144[3453];
	assign cj_6144[5692] = ci_6144[5540];
	assign cj_6144[5693] = ci_6144[2443];
	assign cj_6144[5694] = ci_6144[306];
	assign cj_6144[5695] = ci_6144[5273];
	assign cj_6144[5696] = ci_6144[5056];
	assign cj_6144[5697] = ci_6144[5799];
	assign cj_6144[5698] = ci_6144[1358];
	assign cj_6144[5699] = ci_6144[4021];
	assign cj_6144[5700] = ci_6144[1500];
	assign cj_6144[5701] = ci_6144[6083];
	assign cj_6144[5702] = ci_6144[5482];
	assign cj_6144[5703] = ci_6144[5841];
	assign cj_6144[5704] = ci_6144[1016];
	assign cj_6144[5705] = ci_6144[3295];
	assign cj_6144[5706] = ci_6144[390];
	assign cj_6144[5707] = ci_6144[4589];
	assign cj_6144[5708] = ci_6144[3604];
	assign cj_6144[5709] = ci_6144[3579];
	assign cj_6144[5710] = ci_6144[4514];
	assign cj_6144[5711] = ci_6144[265];
	assign cj_6144[5712] = ci_6144[3120];
	assign cj_6144[5713] = ci_6144[791];
	assign cj_6144[5714] = ci_6144[5566];
	assign cj_6144[5715] = ci_6144[5157];
	assign cj_6144[5716] = ci_6144[5708];
	assign cj_6144[5717] = ci_6144[1075];
	assign cj_6144[5718] = ci_6144[3546];
	assign cj_6144[5719] = ci_6144[833];
	assign cj_6144[5720] = ci_6144[5224];
	assign cj_6144[5721] = ci_6144[4431];
	assign cj_6144[5722] = ci_6144[4598];
	assign cj_6144[5723] = ci_6144[5725];
	assign cj_6144[5724] = ci_6144[1668];
	assign cj_6144[5725] = ci_6144[4715];
	assign cj_6144[5726] = ci_6144[2578];
	assign cj_6144[5727] = ci_6144[1401];
	assign cj_6144[5728] = ci_6144[1184];
	assign cj_6144[5729] = ci_6144[1927];
	assign cj_6144[5730] = ci_6144[3630];
	assign cj_6144[5731] = ci_6144[149];
	assign cj_6144[5732] = ci_6144[3772];
	assign cj_6144[5733] = ci_6144[2211];
	assign cj_6144[5734] = ci_6144[1610];
	assign cj_6144[5735] = ci_6144[1969];
	assign cj_6144[5736] = ci_6144[3288];
	assign cj_6144[5737] = ci_6144[5567];
	assign cj_6144[5738] = ci_6144[2662];
	assign cj_6144[5739] = ci_6144[717];
	assign cj_6144[5740] = ci_6144[5876];
	assign cj_6144[5741] = ci_6144[5851];
	assign cj_6144[5742] = ci_6144[642];
	assign cj_6144[5743] = ci_6144[2537];
	assign cj_6144[5744] = ci_6144[5392];
	assign cj_6144[5745] = ci_6144[3063];
	assign cj_6144[5746] = ci_6144[1694];
	assign cj_6144[5747] = ci_6144[1285];
	assign cj_6144[5748] = ci_6144[1836];
	assign cj_6144[5749] = ci_6144[3347];
	assign cj_6144[5750] = ci_6144[5818];
	assign cj_6144[5751] = ci_6144[3105];
	assign cj_6144[5752] = ci_6144[1352];
	assign cj_6144[5753] = ci_6144[559];
	assign cj_6144[5754] = ci_6144[726];
	assign cj_6144[5755] = ci_6144[1853];
	assign cj_6144[5756] = ci_6144[3940];
	assign cj_6144[5757] = ci_6144[843];
	assign cj_6144[5758] = ci_6144[4850];
	assign cj_6144[5759] = ci_6144[3673];
	assign cj_6144[5760] = ci_6144[3456];
	assign cj_6144[5761] = ci_6144[4199];
	assign cj_6144[5762] = ci_6144[5902];
	assign cj_6144[5763] = ci_6144[2421];
	assign cj_6144[5764] = ci_6144[6044];
	assign cj_6144[5765] = ci_6144[4483];
	assign cj_6144[5766] = ci_6144[3882];
	assign cj_6144[5767] = ci_6144[4241];
	assign cj_6144[5768] = ci_6144[5560];
	assign cj_6144[5769] = ci_6144[1695];
	assign cj_6144[5770] = ci_6144[4934];
	assign cj_6144[5771] = ci_6144[2989];
	assign cj_6144[5772] = ci_6144[2004];
	assign cj_6144[5773] = ci_6144[1979];
	assign cj_6144[5774] = ci_6144[2914];
	assign cj_6144[5775] = ci_6144[4809];
	assign cj_6144[5776] = ci_6144[1520];
	assign cj_6144[5777] = ci_6144[5335];
	assign cj_6144[5778] = ci_6144[3966];
	assign cj_6144[5779] = ci_6144[3557];
	assign cj_6144[5780] = ci_6144[4108];
	assign cj_6144[5781] = ci_6144[5619];
	assign cj_6144[5782] = ci_6144[1946];
	assign cj_6144[5783] = ci_6144[5377];
	assign cj_6144[5784] = ci_6144[3624];
	assign cj_6144[5785] = ci_6144[2831];
	assign cj_6144[5786] = ci_6144[2998];
	assign cj_6144[5787] = ci_6144[4125];
	assign cj_6144[5788] = ci_6144[68];
	assign cj_6144[5789] = ci_6144[3115];
	assign cj_6144[5790] = ci_6144[978];
	assign cj_6144[5791] = ci_6144[5945];
	assign cj_6144[5792] = ci_6144[5728];
	assign cj_6144[5793] = ci_6144[327];
	assign cj_6144[5794] = ci_6144[2030];
	assign cj_6144[5795] = ci_6144[4693];
	assign cj_6144[5796] = ci_6144[2172];
	assign cj_6144[5797] = ci_6144[611];
	assign cj_6144[5798] = ci_6144[10];
	assign cj_6144[5799] = ci_6144[369];
	assign cj_6144[5800] = ci_6144[1688];
	assign cj_6144[5801] = ci_6144[3967];
	assign cj_6144[5802] = ci_6144[1062];
	assign cj_6144[5803] = ci_6144[5261];
	assign cj_6144[5804] = ci_6144[4276];
	assign cj_6144[5805] = ci_6144[4251];
	assign cj_6144[5806] = ci_6144[5186];
	assign cj_6144[5807] = ci_6144[937];
	assign cj_6144[5808] = ci_6144[3792];
	assign cj_6144[5809] = ci_6144[1463];
	assign cj_6144[5810] = ci_6144[94];
	assign cj_6144[5811] = ci_6144[5829];
	assign cj_6144[5812] = ci_6144[236];
	assign cj_6144[5813] = ci_6144[1747];
	assign cj_6144[5814] = ci_6144[4218];
	assign cj_6144[5815] = ci_6144[1505];
	assign cj_6144[5816] = ci_6144[5896];
	assign cj_6144[5817] = ci_6144[5103];
	assign cj_6144[5818] = ci_6144[5270];
	assign cj_6144[5819] = ci_6144[253];
	assign cj_6144[5820] = ci_6144[2340];
	assign cj_6144[5821] = ci_6144[5387];
	assign cj_6144[5822] = ci_6144[3250];
	assign cj_6144[5823] = ci_6144[2073];
	assign cj_6144[5824] = ci_6144[1856];
	assign cj_6144[5825] = ci_6144[2599];
	assign cj_6144[5826] = ci_6144[4302];
	assign cj_6144[5827] = ci_6144[821];
	assign cj_6144[5828] = ci_6144[4444];
	assign cj_6144[5829] = ci_6144[2883];
	assign cj_6144[5830] = ci_6144[2282];
	assign cj_6144[5831] = ci_6144[2641];
	assign cj_6144[5832] = ci_6144[3960];
	assign cj_6144[5833] = ci_6144[95];
	assign cj_6144[5834] = ci_6144[3334];
	assign cj_6144[5835] = ci_6144[1389];
	assign cj_6144[5836] = ci_6144[404];
	assign cj_6144[5837] = ci_6144[379];
	assign cj_6144[5838] = ci_6144[1314];
	assign cj_6144[5839] = ci_6144[3209];
	assign cj_6144[5840] = ci_6144[6064];
	assign cj_6144[5841] = ci_6144[3735];
	assign cj_6144[5842] = ci_6144[2366];
	assign cj_6144[5843] = ci_6144[1957];
	assign cj_6144[5844] = ci_6144[2508];
	assign cj_6144[5845] = ci_6144[4019];
	assign cj_6144[5846] = ci_6144[346];
	assign cj_6144[5847] = ci_6144[3777];
	assign cj_6144[5848] = ci_6144[2024];
	assign cj_6144[5849] = ci_6144[1231];
	assign cj_6144[5850] = ci_6144[1398];
	assign cj_6144[5851] = ci_6144[2525];
	assign cj_6144[5852] = ci_6144[4612];
	assign cj_6144[5853] = ci_6144[1515];
	assign cj_6144[5854] = ci_6144[5522];
	assign cj_6144[5855] = ci_6144[4345];
	assign cj_6144[5856] = ci_6144[4128];
	assign cj_6144[5857] = ci_6144[4871];
	assign cj_6144[5858] = ci_6144[430];
	assign cj_6144[5859] = ci_6144[3093];
	assign cj_6144[5860] = ci_6144[572];
	assign cj_6144[5861] = ci_6144[5155];
	assign cj_6144[5862] = ci_6144[4554];
	assign cj_6144[5863] = ci_6144[4913];
	assign cj_6144[5864] = ci_6144[88];
	assign cj_6144[5865] = ci_6144[2367];
	assign cj_6144[5866] = ci_6144[5606];
	assign cj_6144[5867] = ci_6144[3661];
	assign cj_6144[5868] = ci_6144[2676];
	assign cj_6144[5869] = ci_6144[2651];
	assign cj_6144[5870] = ci_6144[3586];
	assign cj_6144[5871] = ci_6144[5481];
	assign cj_6144[5872] = ci_6144[2192];
	assign cj_6144[5873] = ci_6144[6007];
	assign cj_6144[5874] = ci_6144[4638];
	assign cj_6144[5875] = ci_6144[4229];
	assign cj_6144[5876] = ci_6144[4780];
	assign cj_6144[5877] = ci_6144[147];
	assign cj_6144[5878] = ci_6144[2618];
	assign cj_6144[5879] = ci_6144[6049];
	assign cj_6144[5880] = ci_6144[4296];
	assign cj_6144[5881] = ci_6144[3503];
	assign cj_6144[5882] = ci_6144[3670];
	assign cj_6144[5883] = ci_6144[4797];
	assign cj_6144[5884] = ci_6144[740];
	assign cj_6144[5885] = ci_6144[3787];
	assign cj_6144[5886] = ci_6144[1650];
	assign cj_6144[5887] = ci_6144[473];
	assign cj_6144[5888] = ci_6144[256];
	assign cj_6144[5889] = ci_6144[999];
	assign cj_6144[5890] = ci_6144[2702];
	assign cj_6144[5891] = ci_6144[5365];
	assign cj_6144[5892] = ci_6144[2844];
	assign cj_6144[5893] = ci_6144[1283];
	assign cj_6144[5894] = ci_6144[682];
	assign cj_6144[5895] = ci_6144[1041];
	assign cj_6144[5896] = ci_6144[2360];
	assign cj_6144[5897] = ci_6144[4639];
	assign cj_6144[5898] = ci_6144[1734];
	assign cj_6144[5899] = ci_6144[5933];
	assign cj_6144[5900] = ci_6144[4948];
	assign cj_6144[5901] = ci_6144[4923];
	assign cj_6144[5902] = ci_6144[5858];
	assign cj_6144[5903] = ci_6144[1609];
	assign cj_6144[5904] = ci_6144[4464];
	assign cj_6144[5905] = ci_6144[2135];
	assign cj_6144[5906] = ci_6144[766];
	assign cj_6144[5907] = ci_6144[357];
	assign cj_6144[5908] = ci_6144[908];
	assign cj_6144[5909] = ci_6144[2419];
	assign cj_6144[5910] = ci_6144[4890];
	assign cj_6144[5911] = ci_6144[2177];
	assign cj_6144[5912] = ci_6144[424];
	assign cj_6144[5913] = ci_6144[5775];
	assign cj_6144[5914] = ci_6144[5942];
	assign cj_6144[5915] = ci_6144[925];
	assign cj_6144[5916] = ci_6144[3012];
	assign cj_6144[5917] = ci_6144[6059];
	assign cj_6144[5918] = ci_6144[3922];
	assign cj_6144[5919] = ci_6144[2745];
	assign cj_6144[5920] = ci_6144[2528];
	assign cj_6144[5921] = ci_6144[3271];
	assign cj_6144[5922] = ci_6144[4974];
	assign cj_6144[5923] = ci_6144[1493];
	assign cj_6144[5924] = ci_6144[5116];
	assign cj_6144[5925] = ci_6144[3555];
	assign cj_6144[5926] = ci_6144[2954];
	assign cj_6144[5927] = ci_6144[3313];
	assign cj_6144[5928] = ci_6144[4632];
	assign cj_6144[5929] = ci_6144[767];
	assign cj_6144[5930] = ci_6144[4006];
	assign cj_6144[5931] = ci_6144[2061];
	assign cj_6144[5932] = ci_6144[1076];
	assign cj_6144[5933] = ci_6144[1051];
	assign cj_6144[5934] = ci_6144[1986];
	assign cj_6144[5935] = ci_6144[3881];
	assign cj_6144[5936] = ci_6144[592];
	assign cj_6144[5937] = ci_6144[4407];
	assign cj_6144[5938] = ci_6144[3038];
	assign cj_6144[5939] = ci_6144[2629];
	assign cj_6144[5940] = ci_6144[3180];
	assign cj_6144[5941] = ci_6144[4691];
	assign cj_6144[5942] = ci_6144[1018];
	assign cj_6144[5943] = ci_6144[4449];
	assign cj_6144[5944] = ci_6144[2696];
	assign cj_6144[5945] = ci_6144[1903];
	assign cj_6144[5946] = ci_6144[2070];
	assign cj_6144[5947] = ci_6144[3197];
	assign cj_6144[5948] = ci_6144[5284];
	assign cj_6144[5949] = ci_6144[2187];
	assign cj_6144[5950] = ci_6144[50];
	assign cj_6144[5951] = ci_6144[5017];
	assign cj_6144[5952] = ci_6144[4800];
	assign cj_6144[5953] = ci_6144[5543];
	assign cj_6144[5954] = ci_6144[1102];
	assign cj_6144[5955] = ci_6144[3765];
	assign cj_6144[5956] = ci_6144[1244];
	assign cj_6144[5957] = ci_6144[5827];
	assign cj_6144[5958] = ci_6144[5226];
	assign cj_6144[5959] = ci_6144[5585];
	assign cj_6144[5960] = ci_6144[760];
	assign cj_6144[5961] = ci_6144[3039];
	assign cj_6144[5962] = ci_6144[134];
	assign cj_6144[5963] = ci_6144[4333];
	assign cj_6144[5964] = ci_6144[3348];
	assign cj_6144[5965] = ci_6144[3323];
	assign cj_6144[5966] = ci_6144[4258];
	assign cj_6144[5967] = ci_6144[9];
	assign cj_6144[5968] = ci_6144[2864];
	assign cj_6144[5969] = ci_6144[535];
	assign cj_6144[5970] = ci_6144[5310];
	assign cj_6144[5971] = ci_6144[4901];
	assign cj_6144[5972] = ci_6144[5452];
	assign cj_6144[5973] = ci_6144[819];
	assign cj_6144[5974] = ci_6144[3290];
	assign cj_6144[5975] = ci_6144[577];
	assign cj_6144[5976] = ci_6144[4968];
	assign cj_6144[5977] = ci_6144[4175];
	assign cj_6144[5978] = ci_6144[4342];
	assign cj_6144[5979] = ci_6144[5469];
	assign cj_6144[5980] = ci_6144[1412];
	assign cj_6144[5981] = ci_6144[4459];
	assign cj_6144[5982] = ci_6144[2322];
	assign cj_6144[5983] = ci_6144[1145];
	assign cj_6144[5984] = ci_6144[928];
	assign cj_6144[5985] = ci_6144[1671];
	assign cj_6144[5986] = ci_6144[3374];
	assign cj_6144[5987] = ci_6144[6037];
	assign cj_6144[5988] = ci_6144[3516];
	assign cj_6144[5989] = ci_6144[1955];
	assign cj_6144[5990] = ci_6144[1354];
	assign cj_6144[5991] = ci_6144[1713];
	assign cj_6144[5992] = ci_6144[3032];
	assign cj_6144[5993] = ci_6144[5311];
	assign cj_6144[5994] = ci_6144[2406];
	assign cj_6144[5995] = ci_6144[461];
	assign cj_6144[5996] = ci_6144[5620];
	assign cj_6144[5997] = ci_6144[5595];
	assign cj_6144[5998] = ci_6144[386];
	assign cj_6144[5999] = ci_6144[2281];
	assign cj_6144[6000] = ci_6144[5136];
	assign cj_6144[6001] = ci_6144[2807];
	assign cj_6144[6002] = ci_6144[1438];
	assign cj_6144[6003] = ci_6144[1029];
	assign cj_6144[6004] = ci_6144[1580];
	assign cj_6144[6005] = ci_6144[3091];
	assign cj_6144[6006] = ci_6144[5562];
	assign cj_6144[6007] = ci_6144[2849];
	assign cj_6144[6008] = ci_6144[1096];
	assign cj_6144[6009] = ci_6144[303];
	assign cj_6144[6010] = ci_6144[470];
	assign cj_6144[6011] = ci_6144[1597];
	assign cj_6144[6012] = ci_6144[3684];
	assign cj_6144[6013] = ci_6144[587];
	assign cj_6144[6014] = ci_6144[4594];
	assign cj_6144[6015] = ci_6144[3417];
	assign cj_6144[6016] = ci_6144[3200];
	assign cj_6144[6017] = ci_6144[3943];
	assign cj_6144[6018] = ci_6144[5646];
	assign cj_6144[6019] = ci_6144[2165];
	assign cj_6144[6020] = ci_6144[5788];
	assign cj_6144[6021] = ci_6144[4227];
	assign cj_6144[6022] = ci_6144[3626];
	assign cj_6144[6023] = ci_6144[3985];
	assign cj_6144[6024] = ci_6144[5304];
	assign cj_6144[6025] = ci_6144[1439];
	assign cj_6144[6026] = ci_6144[4678];
	assign cj_6144[6027] = ci_6144[2733];
	assign cj_6144[6028] = ci_6144[1748];
	assign cj_6144[6029] = ci_6144[1723];
	assign cj_6144[6030] = ci_6144[2658];
	assign cj_6144[6031] = ci_6144[4553];
	assign cj_6144[6032] = ci_6144[1264];
	assign cj_6144[6033] = ci_6144[5079];
	assign cj_6144[6034] = ci_6144[3710];
	assign cj_6144[6035] = ci_6144[3301];
	assign cj_6144[6036] = ci_6144[3852];
	assign cj_6144[6037] = ci_6144[5363];
	assign cj_6144[6038] = ci_6144[1690];
	assign cj_6144[6039] = ci_6144[5121];
	assign cj_6144[6040] = ci_6144[3368];
	assign cj_6144[6041] = ci_6144[2575];
	assign cj_6144[6042] = ci_6144[2742];
	assign cj_6144[6043] = ci_6144[3869];
	assign cj_6144[6044] = ci_6144[5956];
	assign cj_6144[6045] = ci_6144[2859];
	assign cj_6144[6046] = ci_6144[722];
	assign cj_6144[6047] = ci_6144[5689];
	assign cj_6144[6048] = ci_6144[5472];
	assign cj_6144[6049] = ci_6144[71];
	assign cj_6144[6050] = ci_6144[1774];
	assign cj_6144[6051] = ci_6144[4437];
	assign cj_6144[6052] = ci_6144[1916];
	assign cj_6144[6053] = ci_6144[355];
	assign cj_6144[6054] = ci_6144[5898];
	assign cj_6144[6055] = ci_6144[113];
	assign cj_6144[6056] = ci_6144[1432];
	assign cj_6144[6057] = ci_6144[3711];
	assign cj_6144[6058] = ci_6144[806];
	assign cj_6144[6059] = ci_6144[5005];
	assign cj_6144[6060] = ci_6144[4020];
	assign cj_6144[6061] = ci_6144[3995];
	assign cj_6144[6062] = ci_6144[4930];
	assign cj_6144[6063] = ci_6144[681];
	assign cj_6144[6064] = ci_6144[3536];
	assign cj_6144[6065] = ci_6144[1207];
	assign cj_6144[6066] = ci_6144[5982];
	assign cj_6144[6067] = ci_6144[5573];
	assign cj_6144[6068] = ci_6144[6124];
	assign cj_6144[6069] = ci_6144[1491];
	assign cj_6144[6070] = ci_6144[3962];
	assign cj_6144[6071] = ci_6144[1249];
	assign cj_6144[6072] = ci_6144[5640];
	assign cj_6144[6073] = ci_6144[4847];
	assign cj_6144[6074] = ci_6144[5014];
	assign cj_6144[6075] = ci_6144[6141];
	assign cj_6144[6076] = ci_6144[2084];
	assign cj_6144[6077] = ci_6144[5131];
	assign cj_6144[6078] = ci_6144[2994];
	assign cj_6144[6079] = ci_6144[1817];
	assign cj_6144[6080] = ci_6144[1600];
	assign cj_6144[6081] = ci_6144[2343];
	assign cj_6144[6082] = ci_6144[4046];
	assign cj_6144[6083] = ci_6144[565];
	assign cj_6144[6084] = ci_6144[4188];
	assign cj_6144[6085] = ci_6144[2627];
	assign cj_6144[6086] = ci_6144[2026];
	assign cj_6144[6087] = ci_6144[2385];
	assign cj_6144[6088] = ci_6144[3704];
	assign cj_6144[6089] = ci_6144[5983];
	assign cj_6144[6090] = ci_6144[3078];
	assign cj_6144[6091] = ci_6144[1133];
	assign cj_6144[6092] = ci_6144[148];
	assign cj_6144[6093] = ci_6144[123];
	assign cj_6144[6094] = ci_6144[1058];
	assign cj_6144[6095] = ci_6144[2953];
	assign cj_6144[6096] = ci_6144[5808];
	assign cj_6144[6097] = ci_6144[3479];
	assign cj_6144[6098] = ci_6144[2110];
	assign cj_6144[6099] = ci_6144[1701];
	assign cj_6144[6100] = ci_6144[2252];
	assign cj_6144[6101] = ci_6144[3763];
	assign cj_6144[6102] = ci_6144[90];
	assign cj_6144[6103] = ci_6144[3521];
	assign cj_6144[6104] = ci_6144[1768];
	assign cj_6144[6105] = ci_6144[975];
	assign cj_6144[6106] = ci_6144[1142];
	assign cj_6144[6107] = ci_6144[2269];
	assign cj_6144[6108] = ci_6144[4356];
	assign cj_6144[6109] = ci_6144[1259];
	assign cj_6144[6110] = ci_6144[5266];
	assign cj_6144[6111] = ci_6144[4089];
	assign cj_6144[6112] = ci_6144[3872];
	assign cj_6144[6113] = ci_6144[4615];
	assign cj_6144[6114] = ci_6144[174];
	assign cj_6144[6115] = ci_6144[2837];
	assign cj_6144[6116] = ci_6144[316];
	assign cj_6144[6117] = ci_6144[4899];
	assign cj_6144[6118] = ci_6144[4298];
	assign cj_6144[6119] = ci_6144[4657];
	assign cj_6144[6120] = ci_6144[5976];
	assign cj_6144[6121] = ci_6144[2111];
	assign cj_6144[6122] = ci_6144[5350];
	assign cj_6144[6123] = ci_6144[3405];
	assign cj_6144[6124] = ci_6144[2420];
	assign cj_6144[6125] = ci_6144[2395];
	assign cj_6144[6126] = ci_6144[3330];
	assign cj_6144[6127] = ci_6144[5225];
	assign cj_6144[6128] = ci_6144[1936];
	assign cj_6144[6129] = ci_6144[5751];
	assign cj_6144[6130] = ci_6144[4382];
	assign cj_6144[6131] = ci_6144[3973];
	assign cj_6144[6132] = ci_6144[4524];
	assign cj_6144[6133] = ci_6144[6035];
	assign cj_6144[6134] = ci_6144[2362];
	assign cj_6144[6135] = ci_6144[5793];
	assign cj_6144[6136] = ci_6144[4040];
	assign cj_6144[6137] = ci_6144[3247];
	assign cj_6144[6138] = ci_6144[3414];
	assign cj_6144[6139] = ci_6144[4541];
	assign cj_6144[6140] = ci_6144[484];
	assign cj_6144[6141] = ci_6144[3531];
	assign cj_6144[6142] = ci_6144[1394];
	assign cj_6144[6143] = ci_6144[217];






endmodule

	`endif